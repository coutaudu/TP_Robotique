��   O�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����DMR_GRP�_T  � �$MA��R_D�ONE  $�OT_MINUS�   	GPyLN8COUNP �T REF>wP�OOtlTpB�CKLSH_SI�GoSEACHMsST>pSPC�
��MOVB RAD�APT_INERzP �FRIC�
_COL_P M�
�GRAV��� HsIS��DSP?��HIFT_ER[RO�  �NA�pMCHY SwARM_PARA#w d7ANGC �M2pCLDE|�CALIB� �DB$GEARz�2� RING���<$1_8k�  �FMS*�t *v M_LIF��u,(8*���M(DSTB0+_0>*_���*#z&~+CL_TIM��PCCOMi�F�Bk M� �MAL�_�EC�S�P�!Q%XO g$PS� �TI����%�"r $DT�Y?R. l*1EN�D14�$1�ACT�1#4V22\93\94�\95\96\6_OVR\6� GA[7�2h7 �2u7�2�7�2�7�2�8oFRMZ\6DE�{DX\6CURL� 
HSZ27Fh1DGu1�DG�1DG�1DG�1DCN�A!1?( �P�L� + ��S�TA23TRQ_Mȫ�/@K"�FSX��JY�JZ�II�JI��JI�D �$U1S�S  ����6Q����+PVIRTUAL3_EQ'� 1 TU_  ��(P���_�_�_�_�_�_ o�_o=o(fVlho�+cAQ�ool�����t<���n���������no�ojo�l�o�o85G�kz�ri ������d��x�)���=L��4�f[�?�\���@�|� ����ŏ׏�����`1�C�U�g�� TU���������:T  2 ����'�9�K�]�o�������<����ϯ ����)�;�M�_�pq�����UP��$$� 1q\�qJ�6�K �J�e��Nm��M͸M����}�Ld�L'�%�L�D�S��E#]`D5�Y޾}Aщ�щ �<�z�9�r�]ϖ�	� �}�ÿտ�����4��X�j� b��u��V߿�������Tnu�Tp��S��� <�N�`��1���� y���������8�J� \��-�������u��� ������4FX )���q��� �0BT%� ��m���/� ,/>/P//!/�/�/�/ i/�/�/�/?���/,? >?P?�/t?�?�?�?i? �?�?�?O�?(O:OLO OpO�O�O�OeO�O�O��O _�O$_6_H_q�,�($1234567890m_U��k_ �_�_�_�_�_�_�_o o)o1oCowogo�o�o �o�o�o�o�o�o+ 7?[�u��� ������)�]��M�i�q��������$�PLCL��ҕ�� DO�?�  ��� 6�O�Z�E�~�i����� ��؟ß��� �2�