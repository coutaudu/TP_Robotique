��  �\�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A9  �����ABSPOS_�GRP_T  �  $PAR�AM  �  �ALRM�_RECOV1�   $ALM�OENB��]OyNiI M_IF1� D $EN�ABLE k L�AST_^  �d�U�K}MA�X� $LDEB�UG@  
����APCOUPLE�D1 $[PP�_PROCES0� � �1��U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $�,NO/PS_SPI_INDE���$DX�SCR�EEN_NAME� �SIG�Nj��&PK�_FI� 	$�THKY�PAN�E7  	$D�UMMY12� ��3�4�GRG�_STR1 � $TIT�$I��1&�$P�$�$5&6&U7&8&9'0'�'�%!'�%5'1�?'1I'1S'1]'2�h"GSBN_CF�G1  8 �$CNV_JNT�_* �DATA_�CMNT�!$F�LAGSL*CH�ECK��AT_�CELLSETU�P  P� H?OME_IO� �%:3MACRO�F2REPRO8�D�RUNCD�i2S�Mp5H UTOBA�CKU0 }�	DEVIC#sTIh�$DFMD�ST�0B 3�$INTERVA�L�DISP_U�NIT��0_DO��6ERR�9FR_�Fa�INGRkES�!Y0Q_�3t4C_WA�4�12J�OFF_� N�3D;EL_HLOG�2�jA�2?�1k@��?�� ���H X�_D�#	 d �$CARD_E�XIST�$FSSB_TYPi�� CHKBD_S�E�5AGN G�� $SLOT_�NUMZ�APREyVD� ��1�_EDIT1
 W� h1G=H0yS?@f%$EP�Y$OPc ~iAETE_OK�B{US�P_CR�A�$�4JVAZ0LACIwY1�R�@k ��1COMMEc@$D�V�QOk@�:Y��G BL*O�U/R , $��1V1AB0~ O�L#eR"2CF�D X $GR� z� S!1$MB_@NFLIC�3\`
�UIREs3��AO}MqWITCHWc/AX_N.0S�=`�_;G0 � 
$WARNM'@0f��@� LI? �a�NST� CORN���1FLTR�eT�RAT@0T�` �0ACC�1�` |�rORI�P�Cxk;RTq0_SF� �!�CHGI1 E[ TT`u3I*p[TY��RpK*>2  x �`� �1�B*HDR�J�* ��q2�v3�v4��v5�v6�v7�v8��v9�PqO�$ <� Mo_oqh�s1�<`O_MOR._ t 0Ev։NG� �0BA � �Qt�Q}��r��@B��v���P�0X����h�`^P@/P�2� �p�JpC_R�bLq�@�J	rL	�$�JV�@�CD�`�m|gv�uMtP_}0sOF� �  @� �RO_����aIT<8C��NOM_�0�1���q3W ���$ !����|hP���mEX�`G�0� �0"�<�`�b
$TFR�J6 �D3��TO�3&@yU=0�� ��YH�2�T1m�E��� �e��f��f���0CPDBGDE���@$`PqU�3�f)����AX 1�dbET;AI�3BUF�F��|���! � ˧��`PI���P�L�MK�MX���[�F>L�SIMQS��wKEE��PAT�`��!� ���}p�C�U� �$}1JB8�`-�}1DEC㺋�p���T� �7P�CHNS_EMP�vr$GA�'��@_xy�q3�`1_FP͔vx�TCR�SPEub�w�q0�cg�S�!�� V`�A���!����JR!0~��SEGFRAp�v r�R�T_LI9N�C��PVF�������Y��P���)B��وD )\�}f�e	�"��	� �.0�Z��Ql�ేSIZCuх�d�T�o�A��ڭ�	�RSINF��p����?�� �ܭ���s���LItx��1��CRC�eFCCC�`��>�R��mR��MAl�R��P� �"$�D�d�c��C��j@TA�����@��l���SEV���jF��_��Fw�N�� ��f��!�� 2���������91C��! ���F�hRG�Ps�
qF���7bg�D���2g�LE	W(��s� �e�>��P�ԒR�D� �&�pou2|��A6�NHANCI�$LG�`-��1�Pd��@�dB�aA?@l���~0R��z�jME��uAk��feRAs3jAZC���T�OEqFCT�q��`F�`m�g�̰�ADI;�  q�� l��`��`�`|��H�S=P�r��AMP��Ĥ�Y8C?�MACES����r�I�$�  *�I���CSX�a�!M�p	$JTpT��X�C_ N�@h�IMG_HEIGH�A��WID��h�VTtE��U�0F_A��8- �@EXP(�cN-%�CU���QU�1w $`TIT�19RISG1ꀿ��?DBPXWO���0= �0$SK���2� DBT% TRN�@ !^�Q0TC�؅ `��DJ�4LAY_CAL�1iR� �'�'PL	3&@�0EAD���'�Q�'�Q�DB��!"�"1�PR� 
� �q�Τ!# T A$�wq$�љL@9$�M?_3Gp� %s?�4Cr�!&�?�4ENE�a�x�'�?_3!0RE\�`�2(H C�p� #$LC$�$@3�B� K��VO�a _D6G�ROS��bcvh�D��AMCRIoGGEReFPAyS|���ETURNcBno�MR_o�TU�`�)�2@EWM��ƒ�GN`��CBLAȍ��EΑ�P��&3$P� 9�'�@�QbU�C�D���0DO�����-DAS�3FGO_oAWAYCBMO����Qme�DCS�C0EVI>@ )3 HJ`1vRBw���gSPIhpJ�SP`wVI_BY��|S�UjHSL�r*XP$��<avVTOFB�\�dFE=A1v�SvTHS�o+ 8�DO?��cnpMC%�d�P��)b�R���  `�?,� $��� J �c #fc ��faסߠebit�cH�fa�"rafWr��dNTV�fbV-pr���؃���g��s?�J�?��0��S�AFE̕v_SV>q�EXCLU�!�����ONL+�<sY��TktOT!!��HI�_V5�PPLY�_,�etw�]fjs_M�8� $VRFY_�#�O�� �v!1��s�bFc"�QG -�0� ~�_��:� 2 `SGn� .�
$����@�A����U�R�EV�-�$��UN��0xK�vU��턍���@��l�i�!q���V�!EFf`I�2/���$FN�X$�OT��@jS$DUMMAY
1ׄ1ׄ�����M�PNIG20 L�����4���A`a�D3AY�e`ADiT� 4��؃5��EF $�
��1�0ѧ�Y�_3�� _RTRQݑ2k D_�Ot@RQ:����'���Y� 21����~�jT|��s�¡3 0��ؑ�	�HגS�U�@��"CAB¡4����$���$ID��PWг�ӕH�g�ViWV_�Ӑ��0�DIAG��q¡5� $$	V�@a�T�ǃ���� ���
0	�R�25��VmE� J�SW��@����(���~���2ZPf~�OH���PP��&�IRs!	�B��7������Aᇀ��BAS9q�z ���iV����4����Cנ�R7QDW�MS9����A�������LIF�E� ����10��N ��
�ɵi���
���^UZi�Cm7QN�@9Y����FLATj�3OV6նHE���OUPPO��w���� _6���d�CT�6 `�pCACHE-�m��Es�B~�SUFFIX��e`� ��@�R�؃6\ԁ2MSW�7bKEYIMAG�C�TM%AH����A��I�NPU��!OC�VIEʠ�!8 �h�� L�d��c?�� 	�!"�9���$HOST� ! R�
0Z�0Z�G�Z�R�>Z�EMAIL\ E��� SBL��UL�G2:"҃�COU���T�DaT�0y�;O $��eSӐv4�IT1cBUFǠ�a�NTf j 5�B��mTC�dA��s#��GSAV<��҅�EK@ b2W�Ppm�PC�e�0ˤ��_��"�`��OTRBu�?P�pM��e���r��Z͓DYSN_�� <��DtU�� �U���T/R_IFS�W�O��A�!=0��/��8��#$@TIKYD#&�L�A����K���/�gDSP��/�PC��IM<���sM�w��Uf�+�XE�p��IP��c/���D  ��T!H0�|�TLA���HS��ABSC$H���F��s�dk�$���oSCi�ʖ�1�!ڤ!>bFUI�DU���c��@PE���C�D�	 ���W�R_�NOAUTO�!?���$���:�PUS�C  �C�"�s�  ��� @H *�LI ��� jUs@�c>
1< 1<G�<R�<��<798999��;�E1R1_1l1�y1�1�1�1�2���GR`�H�l2y2�2�2��2�3�3E3TR_3l3y3�U3�3�3�4����EXTz�NaA <���� �]V� �jU��7��pF�DRi�BT ��	���ò�17ò�REM��FQ̲O�VMb��5A�9TR�OV�9DTG�JMX#LIN�98PJf�'IND2@ʲ
^H* ^s�$DG
�X+��@M`ɵ��D��@R�IV�U̲GEAR�b�IO��K�2ʴN $��HY���_p�`�a̲Z_MCM��ñ�0v,�URwC ,��Wq?  �p?�0P��?0QE0op8Q�aCOԐO`�D��n�P1av�RqI�QTz�UP2�p3E G���TD��os��S0�HQ�W�UNP|SB;AC��F TP���T�Ł)]qG�U%��8� t IFI�� 0XP]`+��UPT̢�q/FMR2�5G���1�s�2LIxaFc�7��O�O�OF��ʵ�2_��N��_������M�F�O�MDGCL�F�DGDYxL	DHQ�D5Ѷ�Oɴ'c�E�HU��i T�sFS��F�I P���xqL`
�s�$EXQ_wq�xwq1��EZ�wq3�{5�v�GR9A�P�4J ��t�SW%�Ot�DEBcUG�#���GR0����UZBKUe O�1  ΰPO�`0��CԐ�t�M�S�`OO��^�SM��`EK�����0_?E K S��P�8P�TERM��L<��*�ORI`��yM��"��SM_�Pd�҅�N����TAǉ�O��$Z �UP>�P� - ��2�K$���L$S�EG�%pELTO���$USED�NFI�<�Pt�� |��
�M$UFR�R���� 6�����`OT���pT���0��NST��PATx���OPTHJI� EH�s� �=�AR��I���8V��<�REL�r�SHFT =���ۘ7_SH:�MO�Ɔ� р��5�O�a�0O#VR��r�&�I��d5U� ^�AY��Q`
��ID�MhS�� q� ERVDx�7 &� h2������!`ӥ�!�`RCXQr�ASY1M"�r�=�WJP�h1�d@EhSב�����U�'�������ђ�P�����V�OR��MF@c�po��tQ�� �U���l�����S�E�_R � h�QTOC6�:�Q��OPbm���*tv�e�1OA�RE���RT�r�O
�]⮒e�R��>����T�e$PWR�@IM0ũ�R_���S�]�w S�P$H�U�[�_ADDR�6H�r�G������vѷR�=p��8�T H�pS ` ���#���#��_���lSEkq�1HS<� �sU $����_Dm0=���+�PR����QHTT���UTH7�V (�� OBJECa!l(Q�Q$�6LE��)_�8�W�px7��GAB__A�Գ�S���I�DBGLV��K�RLp�HITE�B�GD�LO����TEM���%B�g�sSS�@7�HW��C���X��\�IN�CPU�rVISIOR���Di���j���j�l �IOLN���Y} �@C��$SL��$INoPUT_u�$0�b��P�@���SLp��Z������IO^@�F_AS]r[�P$L�P���Q-�.Uƀ)�T��� ���z�HY�7T�-�z��wUOPZu\ `� r�6BBD�B@K���B�P90�����K�����u݀UJ�6] �� �PNEV�JO�Gk���DISBcJ�7/�OF�$J8�	7W IT�'97_LAB���) Q�APHI�`Qt(mDypJ7J���0�p_KEY�`� �Kk��0\s^� �@��V��{6�C�TR퓵FLAG��rLGʴ_ ��9`y8���sLG_SIZ�ԧPXp�FDI"Q� 
��	�� Xp���9����2@SCH_H��R�R� N�r`~���@�p�q��1�`UH�����L#�DAU%EAP�k�ܴ3") �GHݲ&a�BOO>�Rat B3���IT�3g$�`/�RE=C|*SCRN� /��DI.�Sl�=pRG Mb�0�,��'����"���S���W�$�$�'�JGM7MNC�HF�'�FN�6Kn;7PRG99UFG8�W�G8FWDG8HL.~9STPG:VG8`XG8n G8RS�9Ho�c;$�CY��3&�'��p�'IUG�[4�'H��&�� <�N2G+9�PPO�RG�:�%�3P/6OC�$�J8EX#�TUI95Ii�#�B�#�C 3�C70;11���AC�ؙ'1��!NO�FANqA�6��`VAIQ ��CL�a��DCS�_HI	�NR��MRO�SX�aVTSIxWjXSvX�(IGN"��4p81�  `UUDEV4;�U!_BU`���b� _�T�B$EM�[���3A��c� _���e�W�Q`m@19e29e3�9aw��R}Q��d �����{�5���%��IDopX�.�4�=a�&��V�fSTs�R4 Y܀�1��` c$E�fC�k��F��f�fR$�!��e LL�B��p W�)�� �C����P����Yd�$_ f :��V����!�s|��C�g ���C�LDPs���TRQ�LIi � �y�tF�LG�b�p�a�s=QD��w=�LD�u�t�uORG �2�r����8��ç�ҙt0�h �� 	�u�5�t�uS��T�p� s�!���}��RCLMC���<�N�������mpMI�Н�i d�yaR�Q� s�DSTB����` ��!'�A�X��� *�C�EXC#ES�q��MO���j����Xa��N�j��k���_A����A�S��pKʴl� \L��$MB�>�LIw��REQGUIRˢ
��O�ODEBU`B��LSpM�m��4�Z��������ND	!ǰ��an�����DC�B$INeЫ!$�� ����PN���C�P�ST�� o��L�OC|fRI&�|eE�X�A��}a���O�DAQ�p
�$3ON�RMF�@ `��iRrJ@\u�����SUP��
`FX��IGGz! q �s�Rs���RsFRtR��%�cιs��޸s��ΐ<�DAT)Ag*�Eq�E�`t�T�N�Rr tN�+MDK�Ix�)YƎPd��a�H/�"dĸ�<Ue�ANSW�!d�(a�Ad�D&�);���ܔ���s ��CU�"V���p7�RR2���t���Z���A��� d$CALII ��GAQ
�2���RINP0�<$R��SW0ʄH�y�A�BC_�D_J2SqE4��X�_J3s�
m�1SP?�< �	PmԔ�3����������Jy��Մ�V_�O�QIMy���CS�KP�z��:S�J<!��Q�3��3�)�$�_AZ����e�EqL�Q���NTE��"bu����7���%p_N��v����a��4�䛒w��DI{����DHc�����x� c$Vв��a$;1$ZbN`b������yH ��$S v�TqACC�EL�QU�ׁd�I�RC��T?�T<�a�c$PSc��rL������s��z�x�BP{�PATHZ����p���3���f�_@6a$� ��M`C���k�_MG�!$D�D${�"$FW���=�`�@p�k�5D}E^PPABN��ROTSPEE�:a��p)�:aDEF�!�k�$USE)_�SP��CO@S�Y� 6� ��YN� �A� ���{��M�OU!NGO� O9L��INC��,��]D'�=��(�ENCS�#����k�%���IN�bI��>����)�VE"Ӡ2�3_U�b�LOWL�QI@���pi�D,@�����dpir��C���MOS�P�ӔMOܰ����PE�RCH  �OV � �1'|a<#�a��� �a2�m"�,����P��A��%LT��З��ך����&�TR�KE$�bAYLOA ���"�� 1��53-��`S�RTI��K�`MOM�B'���2����\
�3��9b5��DU����S_BC?KLSH_C��5 &D ��°4d�:<+�CLAL`�p��A0���5CHK�p:�eSRTY�@(� �@�e$�<�_�c$'_UM��=ICJC$�SCLWD� LMT��_L6���pE��|GEvM�@�Ku@���E����Ц1
� �Du(PC�B!u(HYp;�(@EC̺�]rXTk�6CNE_%�N�S7V׃S�P� g(V��c|V�Qȟ�{UXC!`HMSH �c%�6l$�{1{�`2���U��$PAGD&;_PFE*3_�pd@�6% �q3)dEJG0xpy�c�OG*Wn2TORQU� ��#� 9l ��"o1l �b_	WY5 4_�e�eT�eI�kI�kI�FE��a��x]�. VECZ�0!��"r1(~pu�<2�/uJRK(|�mr`v��DBL_S�M7��M��_DL�GRV�d�t��t�qH_�S�s����zCOS�{/0�xLNop
�+u����@��aH�6��a�uZ��&�qMY����rT�H�}��THET0�NK23�т��CBֆCB�C  �h����d	��	�ֆ�SB�'��GTS���C��,��S&��P�S�6�`�E�$DU @И��
�G������r]1Q�2�$NE䂗�I�(C�2R���$��ŁAɅ����u�x�qLPH�uВ�ВS'�C�6�C�E�ВT�Pm�W�t���V�V	�T�,�V;�VH�VV�UVd�Vr�V��V��H�-�3�+��QJ�H�UHV�Hd�Hr�H��UH��O�O�O���*�O;�OH�OV�O�d�Or�O��Ot�F�В��R�6�W��SPBALANCE�Զ�ALE>�H_ɅS�P��'���6���E�PFULC���½����E���1uLUTOy_@=eT1T2�V�2N�1q�)�6���@:1�������U1T� �O{�c�`INSE9Gq��REV��ΓDIF�%��1vl����1w� OB���1�sg72x`)�A�t?LCHWAR���AB�Qi5$ME�CH�����(FAX1P�D,����Їx 
-�aO�|ROB% CR�"o�!R�y��MSK_|��9�z P !�_� RV����$1zR�����4�����IN|��MT�COM_Cp=�{�   ��v�$NORE��������| 4�`G�R�b�FLA|�$XYZ_DA��B`��DEBU?� X��$�} ��$�wCOD�1 o��>2�90$BU�FINDX� �^�MOR��~ H��W0e��6��58�4��J�&Q��@TA�� _�g2�G�� � $SIMUL'`v�Xx#�#OBJE��>ADJUS1$ OAY_I>az(DR�OUTG`>�W0_[FI=��T�` �	��I��Ф`� ��в��%D� FRI4�3�T�5ROg`��E�a� �OPWO�np���,|�SY�SBU⠙�$SO!P���1U���PRUN��<PAB��D;�s _m �B1��ABc��@m /IMAG�1�ฐ�P��IM��IN��pd�RGOVR!D�- oPq�xP��L_	ЄQ�<B�WPRBXP���AMOC_ED��� �@�N�M"�A�0MYc19�A��SL������ x $OwVSL[�SDI� DEX@SR&OS�!p"	V�`m%Nw!�aj� �u#�'�(%"Z���_�SET�`��� @0�`�"6�1RI�0�
�&_��'�!�!p���/ lP ���yT�<`ATUS~0$TRC��� ��N/3BTM87"1IY�#$4�A3 ��� �D��EmV",2�E���-1�� �0-1EXE30)A!�2�2f4�#1�� ��20UPI�1s$�ИXNNX7�q#$q[9 �PG��� � $S�UB!16��!!1�#J_MPWAI�PPz#�9ELOy@9���$RCVFAIL#_C��RP<AR�  ��)�QjPATs��E��R�_PL�#DBTB8<anRRPBWD~F�3UMl`�DIGT��<ћ�
BDEFSP>H� � L��3���@_�@7�CUNIr]7�@�1R�0Ҥpk_L��P+1f��	P����k�e`�qЭ J���N��KEQT@R�`W�HPP�B�� hB ARSIZEw�:� I�Q�S/ OR�#FORgMAT��DCO5 ,�Q~�EM%��T#S�UX� �"	�ALI��B��  $>��P_SWI�ЏA�1qp�@�@AL_ �� $�A���B�!��C��DY$mE�1�,`C_�A>� � �@�d���(aJ3r����TWIA4�i5�i6��MOM��c�c�c�c4�c��BP@AD�c�f؝c�f�cPU
�NR �du�cu�b���R���� C$PI ǖoe��od�tWu�sWu �sWu��vm{ �r�[!�P�j!{�$�6�S/PEED��Gb�t QE�D�v�DQE�@� �v���x�A��AQESA�M����Z��w[�QEMOV�򊔉��Л���H�����@1�䶄2��@� ��`��%`�H<���IN�%`>������QB�2�	�2�R�G�AMM~Ʒ�I�$GGET���;D_dz��
1�LIBR�1�GrIT�$HI�0_��;0��ǖE��ԘAΞ��LWɝ����3��[b%�MTN�+aC�E����  $PDCK�$�;_=�� ��$bph $a؅���c���f��)c� �$I� R�"�D�����1rD��L�E����!�[h�>n`MSWFL?�FQ� a�И��Pq�UR_SCR�3`�-��#S_SAVE_�D�~��3NO_`C �!�2`d~���ojXv�� qy��0��ۻN��� �v�̀Ja` <����� ���������x�v�@�|�x�6Û��1o����PM2u� � ��YLQs��؇Pу�@ɣ�Ǟc����W��w�����p����2��M��(�CL'�(a�C&"l�"&�q/!PL�Mo��� � 9$���$W~���NG�ya~�8d|�?d |�Fd|�Md�@��᪐(c�%`X9POGc$a�Z��P@ �� pB ��ʣUv��ҿ������_a_�� |B oi~��i��c��@�c~��j����jE@ F�� �Ü�U��\��z`��P�Q�PM�� QU_� � =8TPQCOU̡^ 7QTH��HO��c�7HYS�PES��b�UEN�t��POd��   ���"U�N40*� 
@O���� P���oE�`�}3GrROGRAG1��2�4O����R����INFO��C ���� ���+q�OI#� (R�SLEQ�vK�uK ��$���D>@����QO�����sƑE�sNU��AUT���COPY���0�j!��M�N� �m��C� �QRGAD�J�ᚓRX�R�$9P.�.W,P�,$�.�s&CEX֖@YC��+qRG�NSD� � ?$ALGOz����NYQ_FREQ���W=��v��T�#L�A��ѫc=��uCcRE�0�#� IF�"���NAc�%�_�G�&3(%���EL�E-@ �jbEN�AB�ҡPEASI _!|���N"�q���&cBՀ��I ����q0f�_`��"AB�!K`�E���pV��'BASUb�%�����0���0$�!6$��� X �" 2� ����@>62=7;QX�ޠR5Pi6*r�-PF��ROGRID�13CB�P��wTY`#�OTO����@��_$!HZ�2C$O ����9��[@PORqC�3\Cv�2SRV )	D6FDI�PT_�p#@�5D��?G3=I"P?G5�=I6=I7=I8!AO$�PF������?$VALU�#q��r$n�FQF��|C [%�����3!�n��PANp�vS0 R�0�Qn�TOeP`���$SPW�I�1:TR�EGEN8ZMROcX�7�s�v���FI�TR�#1B8Q_St��WMP��#Vѵq�U�q<!GRTb�Q�Slì� nSV_H�0DAY��P�PS_Y�����mSo�ARY�2�+0�CONFIG_SE_�PBn�d2��m�8+q���4� 4W�?8�vv[�6�PS~����� @W�MC_F,l�|�a�L�~��SM����a�bNsp����c� ,R�cFL�Г���YN�`�|Mf0C���9PUց�LY�ᦛ�DE�LA4pb�Y��AD�Y�W`QSKI�P�ŧ ľ���O���NT��o1^pP_ ����}w`��ҵ��w�Q �y�Q�yV@�zc@�zp@��z}@�z�@�z�@�z9��q�J2Rf���fbEX��T�C� n�C��0rC���qW`wRDC֩ ���R塘�M�ͅ����f�<��w�RGEA�R� �]��E�D��ڝ�ER��a^�C~UM_�C�p�J2TH2N���4� 1� ���0I�1�� �l(�4�\#����T3PE���DO� ]�����T���O3S���Ւ��~�Xp&�2.�� 4�F�X�j�|����&�3.����ß՟�����4.��.�@�R�Pd�v����5.����@��ϯ����6.��(�:�L�^�p����7.������ɿۿ����8.��"�4�F��X�j�|��SMSK�� 6��'�bP:D�s�EMO& ��f`�6�V4�IIOT�I���P�1��POWER�� �6�pa�Yp&�T ���e��$DSB � �!T/pC�Tb^t�S232:ն� �*�DEVICE�U�". t�RPAR�ITY�.!OPBI�TSFLOW0`T�R�� R+P���RCU���r UXTAS�K�RINx�FAC���1"��ZqRSCHR���b�`_sC����POM�tbPGET_�@�b� g0����P[����� !��$USA@p�1���� O�`�� ��'`���_ON��P����WRK�����D�P���FR�IEND 1x $�UF��#w�TOO�L~�MYH�`t�L�ENGTH_VT��FIRM`���U �E�е�UFINV� �RGI<�MAITI�r���Xzq�� G2 �G�1�1U���+�0_y�|O_�Х���`�#� ����@TCs�8��D� �G߀1#
b`��`�����bo
`�.%�S0#�R ���|����X ��*v0L�T�H�0� �&����)$W�0��EDRpLOCK6'Aqwp�QUi�Q$�20���4�.�R:�1F�5�28�2�38�3F���G��@!�����S���SV�P
��VVV@�`b`���b��so :�|+e p�qP]P�!� ��S��U����A9@�'PR�P�&��S�S�q� �q���2� 0�0�20�haV#�A�����E U�{r
��S��� �c!RXAQ{2$P`N��,`�BHAn�L��r^w2THIC.� p�apC��TFERE)N1t5I�@H.�w1aI8��3��K0G1�(��4���9�r��6_�JFGPR�`}q�b�C� <q� *R� }r�C �-F{� ���ҢA  2�� �Sx����	Od �$��Du���E�C$Pn4�CDSP��FJOG�P�p`_	P�q:�O�1Fu��� nL�KEP��IR�Ad�D]`MUAP&B�E�%P�4�S`��@�R�PG:VBR�K`�5�0n0I���  aR�clR�Br Ax�R�C�@BSOC�F�J�N�UD#`Y15��q$SVDE�_OP9dFSPD�_OVR�a<pC��`�R�COR�W��N����VF�1�V�@OV��ESFjP`c�F�3f�!�CHKh��"L�CH2rFuRECOQV�T���@W"pM�P��e�@RO8�Q�@_�h0a0 @���VsER�p��OFS��CN@��WD�Q�d�Q��Q��U�PTR,�| �#@E_FDOV�MB_CMb�	pB�@BLs"�B+rs!�$�V�	��� ucbG,w?XAM=SpZ mu�b�_MCpE�ހOӞ�`T$CA�@ހD:hR�pHBK��6�qIO8��upсPPA�z��y��u��upҹbDVC_DB��C��1��D��b�!"[�1c��s[�3c��` ă�U��@�QUK�@O�CAB�@7��� Жc� fx
�OzpUX~�6SUBCPUr2�@SQ��sUt��*#��3#Ut���Q$HW_C��D@pH��A.c0�$UNI�TuTo�h�ATT�RI-P|��@CYC=LycNECA��S�FLTR_2_F�I�4�خ����1LPx�K�0�0_SCTvF_h�F_r������FS��Mrm�CHA�Q��<�Lr:�;�RS�D�`�҅Q�3s1p�_TjxPRO��s0�KEM��_�`iST)��:! )�C!��D�I���4RAILAiCQ��Mz@LO�P��T7t� ���!��V�sPRE�S�10��C7���	�cFUsNC�R�"RIN� `s�2�Ġ:�/�RAK�� �pc�p�tc�gWAR�3�pBL|�y���A��������D�AsPd�θ����LD@���P���o1m��!���TI�"�xac0�$��RIA���AF�P�Aä`G�p�[S�ʓMOIs�vDF_��Jc��C@�LMOsFA��HR�DY�ORG��H�]�v2�ְ��MULCSE��-S�L!���J�ZJ�Rg	kFAN_ALMLV,���WRN�HAR�D`в��� ��n�2$SHADOW` �0��AMU_�`�6�AU� R.�F�TO_SBR9��յ@���h�9�B���MPIN�Fa0~�������p��p�`|A�  �d�$!�$��� xBbA}@�� �2SEG���C�P%�#AR�@���U201�ܺ�?UAXE�GRO%B�FW��fQ_t�SCSYrP_�hP��S��GWRI��8�*!G��STR�E��gP�PE"j�K@A�oҽ �B��a���!�P�pO�TO��K@�`AR�Yn3+�䡘�UA�AF�IHP�C$LINQK��~1K�/!_��Ҹa@��!r�XY�Z:�}�5��OFF��`J�r�f�/�B�@/����a��3���FI����:1�R�T/��D_J�AIB�RW���e����S�TB�!��YC��.VDU��b?���TUR�XÒ9��X���pAFL0 g`ǃ2� �����8�R�a 1�JK@K�@M�4?�9��p��"��cORQ���Ai���3H� EP�0����!`-S�ATrOVE|�2M��1�� ��Ӗ�IГO� �j��E4��H��1 }�@�d��1�}�`%��%��AER�A
m�	��E��1@�]$	A!c0��[���7�ձ҆ձAX�cIBձ ��Q�L�%���)���) ���*���*�P�*���*� �*�*1H��&�� �)\0�)\0�)\0�)\0 �)\09\09\0/9\0x?9\1P9DEBU@�$;�Gӯ� A�bn�ABէ�q�Qv[@Ġ�r
Bl�7!CEb�OG �OG��OG��OG�QOG ��OG�OGM�^ G�\���LAB��A<�I�GRO��A@��pB_��D&���S ����F,QB(U��4VAND� ��R$��w�U!��qW �q��v�X0Ʊ�X��v�NT'��}	��SERVE�PN�� $��g�Axa!�PPO�b��px%��Q�S_MRA�_� d ԰T�`�xdERREsC�T)Y.���I�pV��#N2aTOQ�$�Lc�H�$��Ee�T�C� � px ,P�d��_V1^2�!�d��
�d2�k2�f�QW�� q�@@�Q�s$W����fldV�����$���w��"jeOC|Ʊ��  k�COUNT�� ��QHELL_CF}G�� 5 �B_BAScRSMR AB��#�i�QSj��cp1�U%bqU2�z3�z4�z5�z�6�z7�z8�wVqR�OO���pݐu�NL���dAB�S͠dpA[CK,FINpT��4��e���.��_P�UՓC��OU�SP���guܡDr�v��чT�PFWD_KAR�7ac aRE�T��P8G�ܱ��QUEm��� }���A�c�I�/C�Css�ڣ?�v�at�SEMR�	�b���<�.P�TY%�SO�!DD�I1����Cс�'u�_sTM�P"�NRQb��s�Eߐ C$KEYSWITCHڣؽ�D�ڄHE��BE�AT����E5�LE(6b����U��F�����SI�DO_HOM�E�OO�REF]PAR��"����2�CԐO��`qaO�P3@�&�IOCM_�YA��@wHK�� yDp�o�RESUb�ςM����ooFO3RCs�ʳ $�Bu�OM6� � @�
D=Â�U��P4�1�֦�4�3֦4�Y���`NPX_AS�Kr� 0qpADD|{�Z�$SIZa�$VA2P�u��TKIP��۠A���``_�����]��S�C�C2`y�FRIF��pS��˩��i�NFe�
�dp��� xx SIObTE��P�SGLѱTY� &����C��ҰOSTMT��P!����BW}ӴSHO9Wř��SV������ �	aA00vTT�ߠ\��\��\���\�5Z�6Z�7*Z�8Z�9Z�AZ�W� \�ʠ\��A]���\���P_�O0�f�1s�1��U1��1��1��1��U1��1��1��1��U1��1�1�1� G���f����؀ɉ��؀��Q �ش�� ����2���2��2��2�2B�2�V��f�3s�U3��3��3��3��U3��3��3��3��U3��3��3�3�U3�4��4f�4s�U4��4��4��4��U4��4��4��4��U4��4��4�4�U4�5��5f�5s�U5��5��5��5��U5��5��5��5��U5��5��5�5�U5�6��6f�6s�U6��6��6��6��U6��6��6��6��U6��6��6�6�U6�7��7f�7s�U7��7��7��7��U7��7��7��7��U7��7�7�7�m7�d�PVP��wUPDJ�� �`�� {r
�PYSLO>Kr� � #�i� f����S �4RB@U5;���pR@8=F�!ID_Le�h5�HIc:I���PLE1_b��4�$	��&;SA�b� h`�0?E_BLCK���2|���8D_CPU�9 $��9�c3�?�4�"P�]�R �|`
P�Wp�q FALA�S�aKC\AUDRUN�ErAJDrAUD���E�AJD�AUD �TB�C�CJ��Xw -$�ALEN�0�D��@?�RA��Rj� W$PI��F1�A
�42WMp]��C���.�ID� jQ&\T#OR�@>[D�a0S��LACEB�0R�@8c0R6`_MA	�MV8�U]W�QTCV�\�Q]WTn��Z�U�ZСKT��a�U]S�aJA�
t$�Mdg�J��D�LU9a]U�A2A�<��`�RaKS"PJKefVK��wa�wa3icJ0l�d{cJJ�cJJ�cAAL{c�`�c�`�fe4�e5�B�QN1�\P�`�[�P.TL'P_���A��@Is� `�0GROUN0�g�}B��NFLICa��=pREQUIRE
�EBUJ��AfY��P2�X��@]v�A��G�� \m�APKPRipCT��P
��;EN�xCLO��y�S_M����yLU
��AL�� �7�M�C�R�P�B�_MG���CF��0$�␉P�%�BRK#�NOL�S�%�2�Rc�_LI�%�i�S��Jr�e�P �diP�ciP�ciP�ciPD�ciP6��߱��8B�����A�t�� fr�B�A ��A�PATH
�#��#���H�N�xp�`CN��CAt�i��r�I�N�BUC-P1y�C�PUM��YPl���l1E�@���@���`o��PAYLOAa�J{2L� R_ANx��LG@��ߙ��$��R_F2LSHR��%�LO�x�)���|7���ACRL_� v�i�r�ה�BHA0�R�$H$���FLE�X�s�AJ�E� :�O�F]Pȧߤ��O�A]P�O�O\F1 ߡ-�A�_)_;_M___q_q�E{_�_�_�_�_ �_�_�_oH�e�g$c edU�w�,o>oPoޡWj	T��F�Xl�bce�� ��ne��zo�o�o�` �e�e�e�e�o�o�oy�rJ!t� � `-?Q��� ATZ�leq`ELȰ *�jlxJS��spJEP�gCTRr�U�TNv��F(�]wHAND_�VB���M0�� $��F2$��sb��<2SW�2��v��� $$M��R >���O������厂��Ao0ܐ�n1$��A(.�10@�AN�A]�/�/��0@�DN�D]�P2=�G]@��STB���4O���N`�DYt@�p $��7��}��ߡ��:�ޗeg�����d�P ������Å̅Յޅ�:�J�u� �ത���"��q�!ASYIMM��fpM��`8h�:�m�_SHrw� ��{��蛟����џ�Jꜛ������.g�_VI����s>	 V_UNI/�$?�'�Jfe6"d6":� :$Q�G$k&Z�`m����|����%������Sdq�pHH@�rݙ�f�!EN��
�DI]���O4`�@� !s�� O�>�I!A ��Q�819@�3F3�08���@;A�1� � ��ME����a2�"�1T� PTq��8��1pt�p��8�1�9T�q $�DUMMY1G�o$PS_X�RF�ֽ�$�6!ALA�#pYP���2�3$GLB_T��5E��01�@��Y�'1� �X�p]w�ST���spSBRM�M21�_VbT$SV_�ER�OWp_CwCC)L3@_BAɰO;2� �GL  EW$q� �4+p�1$Y�ZB�W�C[`$���Ab0肒��AU�E� ��N�@v0E$GIni�}$�A �@8�C�@$q� L+p�F�r}$FrWNE+AR��N_�FLY���TANC_���JsOG?��� ��$JOINT�!xq�1�AMSET$q��  �I3Tʱ��SpM�U��$q�����MOU��?�spL?OCK_FO9����0BGLV\�GL��XTEST_XM��p�QEMP�P��xb1B�P$US~1��@� 2�sp�C@a��b���P@a�aACE�pSa` $KAR��M3TPDRA8�@~duQVEC�f�yPIU@a�EaHE��PTOOL!��cVv �RE�`IS3�r�d6ÁU�ACH�P�S���aO[��3�42��PSI�r � @$RAIL_�BOXE�!spR�OBOd?�aAHOWWAR��0q�0�aROLM�2Vu�р�dgr��p�T�a���^�EOU�R� H R^cI2���P_$PIPfN����br�ag�@a�p�P���OH0 � D�pGLOBA�6��P����3@�r8�S;YS�ADR7�� �0TCH�� � ,��EN�"1A
�Q_�Dp����R�VWVAd1� Ǥ �`�B5PR�EV_RTq$�EDIT��VSHWR��KFԀ���A��Ds0
���H�EAD�� ��潃KE�A�0CPS�PD�JMP_�Ld 5��R��#4��Ue�I`S7�C}��NE�`8�s�TIC�K!�+M5�F�H=NAA� @�pc���$�_GP��v&@gSTYj��aLO3A�qQE������ tk 
��Gv�%$����D=K@S�!$@,!� x1E50FP��SQUx`�B��TERC�0��TS��� �&AW@�� ����x��aT�O�0�3Fc�IZD�AE�1PROC�2Ѣ1�psPU#!�_DOQR�o�XS�PK 6AXiI �zsEaUR��ɳ8�7p��.����_,�`@�ETA�P�R�����F�
t�R~���l �� ��ꔵ�榹�� �� ���0�ڵR�ڵb� ڵr��͟��*��
��s��C)�k}�����SSC@ o� h�@DS���1�0SP20�AT�`��⡠�o��2A_DDRES�cB���SHIF��7`_2+CH7�*�I:@X���TXSCREE�����TIN!A�CPk��D�qB��C@� TU�z@Ţ 8�yAV@���7������RRO; fP7��ر�W4�qUE$4� ��� Y��0S�A8�R�SM���UNEX0k� 6"�� S_�CB�@%2�E�`�%B�C�R��� 1�t�U�E{��,2�B��ѠG+MT~ L�!�f@�O�v�$$CLA~<� ������ՠ�p����VIRTqU� ����ABS�����1 ��� < ��;�M�_�q����� ����������% 7I[m��� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?^;���GAXL��B���+�7  �p4INy?�1�o4��_EXE�8�0�6_UP�м1#����LARM"�O�V ��2l4L�M_P���d^?BOTO fOxO�J0O�O�O�O�O�M, 
6�_j6�NGTOL  �#�	 A   �L_^[�PPLICf��?��0�P�Handl�ingTool ��U 
V8.1�0P/11  ~S-C�(
ya�SW�RՠԄ�Q
F0�Q�U����ՠ
1232��TOh��X��Z��`��7DC�1�P\�SNone�  EL@T�FRA_ 4��YWbl�PpQ��TI�V�5�S�3�cUTEO�� A�4�9P1�GAPON��n���`OUPL�p1I� �`&tg9�`UB� 1K) ��0x0|0|�p���s�1�s����� ��Uvt�H_ur�zHTTHKY���cu� ���#�}�G�Y�k� ��������ŏ׏��� ��y�C�U�g����� ������ӟ���	�� u�?�Q�c��������� ��ϯ����q�;� M�_�}���������˿ ݿ���m�7�I�[� y�ϑϣϵ������� ���i�3�E�W�u�{� �ߟ߱���������� e�/�A�S�q�w��� ����������a�+� =�O�m�s��������� ������]'9K io������ ��Y#5Gek��|BuTO6P�o�cDO_CLEAN�o|@t#NM  ;[_Q/c/u/�/�/4�_DSPDRYRL/?uHI�`/-@@/ ??+?=?O?a?s?�?��?�?�?�?�?<xMA�XrP����g�1X���Q�b�Q�bPLU�GG�`��c�ePRUC� B- �+�/��?WBO\B�/@tSEGF�`K�O�G�A-/ ?/__+_=_O_�O�ALAP�/�N�s�_�_ �_�_�_�_o!o3oEo�Woio{o�cTOTA�LFHI�cUSENU�@�k ��o��BpRG_STRI�NG 1�k
��M�`S}j�
q_ITEM1v  n}m6HZ l~������ �� �2�D�V�h�z����I/O S�IGNALu�Tryout M�odeuInp�̀Simulat{edqOutތOVERR� � = 100rIn cycl҅�qProg A�bor�qȄS�tatuss	H�eartbeat�wMH Fauyl\�e�Alero� ��������ß՟���8��/� �{ �(2���������ȯ گ����"�4�F�X��j�|�������ĿF�WOR�@{��p�ֿ$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D�8V�h�z�PO{P� ��ˉ���������� �/�A�S�e�w��� �������������DEV��D��1�k� }��������������� 1CUgy�����PALT \����"4F Xj|����� ��//0/B/T/�GRI@{�! f/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?z/�`R\�0A �/
OXOjO|O�O�O�O �O�O�O�O__0_B_�T_f_x_�_�_OPREG��PHO�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
.�@���$ARG_���D ?	�����q� � 	$��	+[�x]�w����y�vpSBN_CON?FIG �{ց�Ղ�qCII_SAVE  ����q�rvpTCEL�LSETUP ��z%  OME�_IO����%M�OV_H9�L�R�R�EP3L��pvUTOoBACK$��}�FRA:\��[ ���V�'�`:��W� {� �� �x �]>�P�}�t��������������� )�;��UΟg�y����� ����L����	��-� ?�Q�ܯu��������� ϿZ����)�;�M�_�>A��dωϛϭ�p�����ϲ�INI� ��T�u��MESSAG����p>�ODE_D>���͆9�OF�H߶�PA�US��!��{ ((O�r�߲ۜ� ����������*�,� >�t�b������{�~��TSK  ��x��Ϲ�UPDT?���d5�U�XSCRDCFG 1�v_������|��������� �����e�0BT fx����������rs��G�ROUN)�i�UU�P_NAf��{	���R_ED�1�
L�� 
 �%�-BCKEDTA-Cz���[��t�]�-����Z�r�W��r/  ���_%2h/y�F/�/<"� �t%�/�/C/U/�/y/a#34?�/�?�/�.]?@�??!?�?E?a#4 O p?MO�?�.)O�O�?�?�OOa#5�O<O_`O �.�O`_�O�OO_�Oa#6�__�_,_�.�_,o s_�_o�_a#7do�_ �o�_�.�o�o?oQo�o�uoa#80�}h �-Y��Aa#!9�lI�4��-%��������a!CR g/�o�&��m�Z���೏I�׏U�NO_�DELasGE_�UNUSE_qL�AL_OUT ���>#tWD_A�BOR��T�I�TR_RTN׀<l�NONS���.�1�CE_RIWA_I)�5�y��FF���.���_PARAMG�P 1�����?
��.��CWp  O��Q��Q�U�Q��Q��Q��Q�U�Q��Q��Q��Q���Q��Q��  DF DI�p����y��ͅ�둴� DU��Ѱ��"Ѱ�*��1Ѱ9��@��.?�y�HE��O�NFIG#���G_�PRI 1�� �Ё$��S�e�wωϛϸ�Ͽ���CHK��19�5� ,5�� �%�7�I�[�m�ߑ� �ߵ����������!�(3�E���OF��찫�tCO_MORG_RP 2֬ h�<���� 	 ���� ����������̣������q?����p��`�:Kh�:��P�a��!��aÃ-��������.
 ��
��r�@�����.�`MCPD�Bc��$  )�cpmidbg0N�� �:�� x��瓆p�������K��
�-���� w�v��j�Igf�� ;f�/��/� mc:,/T/~kDEF "(ր)@ cebuf.txt`/�a/�}�_MC��u� ԰ d�%�#����-���!5Cz � BH�B����B�H'B�`�C�B�r-�CZ���D�36C�G�C���D@OC���kD�w�Z=E���E�OE���\E�dE��	F��	�� ;��"4���S<	j��4~j��������A�x���C\Q�DD�i�D@Z>N@ �DE�D�  F��E�oF`[/R�> �JBEL@�Gb��FO�\�G�L��:�  �>�33 ����;  n��;�#5Y�E��; Aa��=L��<#�
�E�O/�"RS�MOFST �.���)T1��DE� �� ��
,�Aj�;��B�O�O^�.TESTy"._�v�R��g��_%6C�4�@���� A��A62��;0Bl�;0C�(@@c��j�:d[�
�QI_���]��QT��FPROG %,���o�UT_IܑZ@䖏��d�KEY_TBL � 6��
A� �	
��� !"#$�%&'()*+,�-./01234�56789:;<=>?@ABCy �GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~����������������������������������������������������������������������������q���������������������������������������������������������������z`L�|��kp�z`ݐSTA�"��T_AUT��O�e��V>�INDTO_ENB+���ROQI�;�T2��t�a�n�v��XCˣ 2�j���8
SONY? XC-56�_	B}�u��@��Ͷ4( А��HR50
���+�y7=�O�Aff[��o��ß �����՟ �0��T�f�A������w���ү�����f,T{RL|`LETE��� w�T_SCR�EEN ,�_kcsc��U���MMENU 1u <*�o�� �������ǿ�&� ���\�3�Eϒ�i�{� ���ϱ��������F� �/�Uߎ�e�w��ߛ� ��������	�B��+� x�O�a������� ����,���b�9�K� q������������� ����%^5G�k }������ H1~Ug�� �����2/	//�A/z/Q/c/�/�)k�_?MANUALÏF��DBCOe�RIG�4�5�DBNUML+IM��:�d�UY`�DBPXWORK 1 fk�_[?m?�?�?�?�]DBTB�_)� !�_�Q��PK4�!_AWAYz�#:�GCP �R9=|P�6_AL0-���2�"Y6��P�(_�DBG 1"ZY�I�,�K?�O�SrO�O��8_Md�I)PL@|+`�CONTIM3����T��F?I
��eTCMOTNEN�D�oSDRECOR�D 1(fk �<�O�SG�O�Qm_ �[B�_�_�_�_xX�_ o_4o�_Xojo|oo )o�o!o�oEo�o 0�oT�ox�o�� ��A�e��>� P�b�t�������+� �������:���E� ͏��������'�ܟK� ՟o�$�6�H�Z�ɟ~��i�w����@eser�ved for Tool ������m�"���X��@mm�y $0E0u� #33Y������ƿ𱿿����@	! T�P Key2 (ABOR�@$�6�H�`��l�ۿe��� Pq�5u�9 گ����X����ώ�C��At Release)q��8u�E�|ߎ����JTOLERENC DsB�IB@L��� �CSS_DEVI�CE 1)�9  �6��)�;� M�_�q�����C��_LS 1*���� �����!�3�E�W������PARAM �+`Ii����_C�FG ,`Ki�d�MC:\��L�%04d.CSV$h�� c��i�A��+CH z� �Oi�Q���'�2�!~|l@0�JPѦ��RC_OUT �-�;m@k���SG�N .�5?R���\�30-M�AR-22 09�:08��?11}4�14:45���� Tnu��-)i�*�o���Im��P�uG��=��VERSI�ON �
�V3.1.j�� E�FLOGIC 1�/�; 	�(�@0����PROG_ENB!OFR�WULS�G �6��_ACC6(A��.C�7#WRST�JN�@�&?R�#DE�MO,(A0E{!IN�I� 0�:�5?1 �v&OPT_SL �?	�&�"
 	�R575i�� 7U4�)6�(7�'5j�
2182�$�6?�>�$TO  �-@t�?�V� DEXd'�d?U�3PATHw A�
A\�?��?O�KIAG_G�RP 25���� �	 E� � F,D FAD�`QC��@IC@��nO�LkA��ЗO�NCe�ECl^OCk�I$C��C�� B�m�I�f362 67�89012345��B�'  �cP�A���A�=q�A�A�33�A�z�A���A��RA���;A�P���JPj!@\@p	 GQ���A�������B4�L��D�(j!
R�P�{A�P��P؜P�P�G��Aď\A��A�Q�*?_Q_cTP�*�б)�^�PϸPU�P� P��P��P���A�ffA�P#P�_�_�_�_o��X_�PZ@`U�PO��
AJPDP>*$P8P2@`,�lWo�io{o�o�]`��A�[�PV�PPPK
=AE�A?P�8��A2�P+ׁ
�o�o�o�X���`�$PLpxPq�Pj$Pc P\Q�;ATPL��bt ����TC@R�Q3a�aKq�p^M=�G��z�>8Q솅^M8���b��7�Ŭ���^M@ʏ\ʆ��p�օE@[PAh�	 �C@<�C�<��t�=�P=�hs=���P�^M;��
.�<#�8�[ �?+���C�  <(��U� 4Ƃ�̝�r����~���@
"?fE6���8���� ��9�k��0�ʟ@�f��H�����~�?Tzᐾ�;�ʥ^M�{��G��^NcQ����^Nx`��7��C��O
�@��CkJ=C���Ck�^M�m����|��ఱ`K
�׿%�ED � E�� ��D+�	�C��O7�j!�8��6з��5���lV�?�6�2 e.2�߫2!��R��M����~Q�C^�������#Ϡ���Ϣ{�����I ACT_CONFI���6������eg� ASTBF/_TTSd'
)B��C#��U���MAqU^ /��MSW���7��_P��OCVI�EWi�8��	 �������*�<� N�I��~������ ��g���� �2�D�V� ��z������������� u�
.@Rd�� ������q *<N`r� �����/&/`8/J/\/n/��RC��	9�5v�!
/|.�/�/��/�/�/#??G?[�S�BL_FAULT� :�*��a1GPGMSK�7t7�0T"A� ;ٵ���MC: �C�O�:|#P��OO1OCOUO gOyO�O�O�O�O�O�O��O	__-_L� �<���1RECP�?�:
�3�_���?�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�oI_���UMP_OPT�IONK�m>qTR��L�q9;uPME|J�.Y_TEM��È�3BK�r�p��ytUNI���MՏq��YN_BR�K <��y8EMGDI_STA�u؂��q�uNC�s1=�� ��o'��|,d�_m��������Ǐ ُ����!�3�E�W� i�{�������ß՟|+ ������[�&�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ���2�  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� �������*�<�N� `�r��������� ����&�8�J�\�n� ���������������� "4FXj|� ������ 0BTfx���� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?��?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_�?f_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<r_ `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�XF�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү���,��,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/� �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObO�/�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6olOFolo~o �o�o�o�o�o�o�o  2DVhz�� �����
��Ro @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ��8�&�8�J�\�n� ��������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ���� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�t߆ߘߪ߼�� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv����� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?� �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_x?f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�oL_&L^ p�������  ��$�6�H�Z�l�~� ������Ə؏���2  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶�������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x����� ����������,�>� P�b�t����������� ����(:L^ p�������  $6HZl~ �������/  /2/D/V/�f/�/�/ �/�/�/�/�/
??.? @?R?d?v?�?�?�?�?��?�?�?I�$EN�ETMODE 1�>r%�     4@�4@<E7OIH@RR�OR_PROG %#J%�LH�OLF�dETABLE  #K|/�O�O�OJ�RRSEV_NU�M 2B  ��-A)PdA_AU�TO_ENB  qPE+CaD_NO>Q� ?#KEA(R�  *��P��P��P��P4P+�P�_�_�_ZTHIS%SLA+@�S[_ALM 1@.#K �LD�\�@+�_;oMo_oqo�o�o�__R`P  �#KQFB�j@TC�P_VER !�#J!�O�o$EXTLOG_REQ�Vs�QY,sSIZ5�'tSTKRyoU��)rTOL  �LADz�R�A 't_BWD�`�pHVܻqDw_DI�q Ar%STDDLAKB�vSTEP��@>�pOP_DOtbA�FDR_GRP s1B#INQd 	�o�r�F@c��[���w��#/�[�7u���� ������c���ɍc�C���Bf��B�[
�A���A�wt�A��aΎ�I�B5YBp�_�@���A��AZ�΍ɏ?�*��c�N���r�����  �A��A�1\�>�����D@
 IJa^�֑Β�׀%�b��ׄE�ݐF,D :�D��`E���)�D  �E�� b�D+��m�C�(�C��N���B�ƈ��΍@7UUU��UU��ۯ�&�8��� E�@����΍OHcG�P)�K��^6�Jk�΍?��R��:G:�z�9�{����΍������>��y�eLA�§�����G�KFEATU�RE Cr%�p�JAHand�lingTool� � svde�English� Diction�ary��
! 4D St��ard�  ff�s��AA Vis�� Master���� R597�n�alog I/O~(�  90 HS��gle Shif�t(�R6417�u�to Softw�are Upda�te  4 RR���matic B�ackupe�49����ground� EditI�  �oadiCa/mera[�F_�4��t��nrRndI�m���duc��o�mm@�calibw UI�� ERm��Con��@�oni�tor��ct\j�3�tr�Reli�abt���PCVL�Data A�cqu=�:���.s�vk�iagno�s��X���cflx�k�ocument�;�eweE���'�O�k�ual Che�ck Safet}y%� g H5���hanced U�s��Fr���PC���xt. DIO� 5�fi�� de�f.��end��ErrD�L������"��s-����rV���� �p��41m�FCTN Menu�йv`���H55��F�TP InF�fa�cv�  J�J�G��pB�k Ex�c��g�� Par��T��Proxy� Sv��  j6�16�igh-S�pe��Ski� �6.fd㰎��m�munic��on1s������urm�F�~_� R67\����connect� 2��04��In;cr��str�z��FCB��KARE�L Cmd. L���ua��J�Uc�R�un-Ti��En�v#�"
c�P�e�l +��s��S/�W��  �License����փ�$�Book(�SyE�m)��! �toMACR7Os,��/O3�{��IF��H���
� 81 ��Mec_hStop��t:��z� T "j�Mi��w� ����Mix���X����orch���odu�witcIh(���o:҉�.� d -��Op;tm� R7*����fil��Pic�k�X�g� OA�D�ulti-T�������v
E�PCM fun�T�z�90#ow�RgegiE��  d���PH�t F* �D/�[Y�Num �Sel6  ry���y�� Adju�����k�w�  {pr�tatuR�*�NDI��ٵ�r���RDM Rob�ot�scove��*�Rem4 �n�� ,���	#Ser�vo� ��?SN�PX b��(�rty �w�LibrÎ��pbo��w�� �E{   m� W oz��tm�ssag� Pv��!z�[s in VC&,Ӧ���` ���(TP6�"/I�� )��� �MILIB=fx�tp� P Fir�m��)�d���n�A�cc����e�71T�X��L��� el	n <I0� �����e\mc�1rq}uu�imulaCѾ�� te.f�1uf� Pa���Ma���T��^Ѡ&��ev�.�Ѧ�USB pYoo @�iP�a��� ��,@nexc�ept��# n�� ��\@�����n0V�C!�r���:hk �1<�j4<�{+�4<�SP CSUI��к��IXC�&roؾHx�� 
�?Web Pl���C97��QC!�Nl2 1R���ԩ�D��3%F�y i�gXGrid!?play o�gXh� ��L� �iRnI/VMRe  e� �-2000iB/�165��rAsc�ii���1�� 5w (K�UUpl��H�35�s!��!t�w rc��Cyct����]ori��5%F�RL��amY*�H�MI Dev�� 1(Y!����PC��-@|o #asswo&��2
49\��64MB DRA�!	�l2��bFRO�kY�7�r�c�visD���5�c���ell[�L�H�54�sh*q�"�0C|c�^�2@Eu���p�6JDEutyt�sH��VIct�� .��� ��sp �2��aV�B by� 
 ��	 B"X�q git2���T1>�nK%.10�OL�`GSupB�Rc�OOPT ��njNS r�bS�B�cro��c	#{%�T mjp���='�a�puest�*�SS�`e�te�x{� ���$LimipYb�Sp����1��0P���gJ�n�Virt��	#����Mdpn�8��h5�1>CVIS� I�RpvC�JDIRC�ALv>D�+�IC�:;0x ��ph�icD�hо�Abuii�l�� FN�!PMM�p�� !�flowh1f.s�k�OSFILE �Ar" u�co g{tp��BMON���IX c�җ!m |T�N@PTTB:��=i��R805� ��J����
��⊔j��^�m����"PA�LT:�`clud����AIW�- Woait/Y�ea�� tk��TP�bD�OES NOT ?RESTO �60�Lin��mark��useJ�z ���c�  Synch�r@�z���DSUP�PR��PRG I�N AR�A ��A�g��OVC_VA�LUE�OBLEkM ��V��TMi�TMW��G���ab��A MOTIO�N�STRUCT� l��BRAK�E ABNORM�x� ��g�$FM�S_GRV0ISM�ATCH=uu�Z�M�AST HANG� UP 37m�M�ULTI WIN�/LOCB���SE�RVO��AG G�AR*�
�GRID� DETECT BUA���!0�����TRANSLAY�?OF UTX���F DB/s�DO PULSE@�ENCCAMER�Aǁ�c�`REMARK FOR�4� w�L�0\h����EXPANDED POS>���%�'����SCREE�l�AY CRUS�H �P!�OTN�560����fԡ�N�D�SYRUNN�I��Ɛ�USR���F TOLp�N�CE ��vK�FS�E��Ŧ ���S-�144 A��AR�T��
p�FA_� �CPMO-073��wAUIs�0��m�pl����ڢ�p!sᇡ�����R��sydem�ַ���A��snosv.�����޷�i���gAQ S���HQ��a_�cmC�-PH�T���!  ORsP�A&;6�`�PR䏡[qdp�(Co(��Y�P,�" �1�Ҁ���G���ҷ�g�R�556�ִ���ic���e�|��G��tg���2�G���aHP spotplugN�sSp��O�-inb�_SPPG ��0~�r�(SC�P`��L8C���J�\sw'���  �� �t���^� ���trsv\<���1.pc
���.  fx_�2�����%3��B	4.:�B��5���"&6�#�C7�	��bB	8���Btn
�P0���=�F�n��sN��Nomi�p Po�si�Q���NN�549~�Ї�`�(B�ѝ���TXP�5
n��os\nm�tp "NMTX" #1�П]�set6�OMP��.����-fxui=fN�-fle��b�FXUFd�Ё�*"�('�6	"$  fC "*!�sq&_�� �o$�	 ,]�t#�w��rl�o(uf�.vr.��'
�@in�cus. ��3&#2+1��"��M? U4K?]?�?�?�?�?�? �?�?�?�?O#OPOGO YO�O}O�O�O�O�O�O �O�O__L_C_U_�_ y_�_�_�_�_�_�_�_ ooHo?oQo~ouo�o �o�o�o�o�o�o D;Mzq���t����� ���	 �  7j$�܎�v|��r�q�j847\wti�v��/���a��/�q���weW ��=����47,r768nR�asyArm&�Gfun?�f�C�R� S01h��Ь�(X�t E����X'��~�\popup�ct�#Ã,��a�N�M�-Shel=ld�R533R��^J� (Mu��-[����;'���vrd�bc2
5C�%� �e�nio.fC�En�H�ced I/ODd��3���J�6v��ŗp��ܷ���rep�a��c���?�acc�uairR�AP�A#irS�6;�0�kz� (\�p���O���S�ca
���4�O� ��2�!S�� 2 G�uc�����49 R#63z����(�����@��g�aΠi1b�#A�oSEL�^�@/���!C�`�n,�aflowL�3� �AF-AS-FM�S�mmP�AFS	M�x�2~勁����(غ����S�˴��afgl
2��G˾!���̴ۢF�̳2V�F�e�AFް���� �����᳣�O/�e�2ȡ̱��d�̱�2L�AF2�Ͻ�2 �����l��RӋ1�B�sŚ���x���!w�����G�_�ɶ3��A8�!㹽�AS ��~� 5������`#����v�LO��.���˱��ݻ��C�clrp�thR�ic C�l[���thϜ77�8��7��gv�ȀBas��@����� �ရ���>�S��㒐��t�pe=���s�sub������n��=�� /�w�set�����"�q��w�q�Off-line Sv�ulari6�>�8�5>���[�85 (� ��tya���si�ad\tp� "SIAD�/�����,k�plug���Dispens�e P� j�=�SPKLG. 9s�(���g-i��� ����ea�\sldsApi�"�U8���0�� L% Trk F ��̀<��>��ꖇ�%���For��t�q���(�]tcyc "T�����k��tgtp�/��!l��la��-#ptkmisc5#�"!�����w� ~��o�sable EOAT<�_�G���� �(@��
� ��3Q!b��"���%1��Fou���os1�)t�47�
���47 (U4��on�)0�_�K1 �2+3��7��a�J5���r70��ervo� Tip Dres�08>���0ȁH7�r7��A?\turnd @b����D�'�����MHb<+�2	��@_��Lq�32]?C5/�S���Ain`�� ���'g�cht ��VG��r~�SGCH J*!�J643>�Q��G�N CfQ��cT\�svsvch��C�H/���Tglgo9uV/�[gnc]����_�P�R�	dV;�sg�dia�Ssb cgorey2XDG�PC70�P�Q{<�b(~d�7�`O��rc�cini�b���^btdw�j95m2Ҵut@unSsCS<���R Jp�iH8r({��u��0��q�Pat݂c��w�����ux�h�869I�7�l;�

/F,
1v���3� mtsv �"MTSV�X�j983\R���&P�s�ov��&_p���/vruk%_c6�p� ����pex_�r�col$Q����Bv�v"�r���&�sxc?M.Tool��xk��=MTOF7p�84 J571 R814�!7E�ǈ��(��q���	mtofs�0��ߘ�2��⒑�pt�a��ll�eto���k�PTLeC�9����J9�813���H���T��4�9��`k{;��1�a\�pmk920 "K���S!R����1�(Ȥ<���2¢2�_�ި4���!�ڣ�a6�1¡4��0����PE�ܣ�q8�4f�4C�c&0�5f�����ݤ���9�7f�7C��ަg�r@"GRIP"�.�쿶��1i "O�PTIC��1ݧpa�lf "PALF��Q��@�{ĻPSS�UC�F!ަcpt "�UNIT�S7mަx=f�XFER��ԃ��et��L�U�&���ŏ��psysd�j��/����mޤopti��Kޥ����7���ssu��+�ޤcpG!W���er��S�N�t�ߞ�sӸ��d+�[��adpՂzaAdapt CtrlF�&3q50E�G0汫���_���l\apa���.�C����a�1l�"�gui� GUI��T���c[�c�l�xogJoU �etra�&��u̞��86F�� (Č��r6��re��3�ETN;���SЗX��5x��j�722\cust�_wv6�RS�v!7x�RS�[8�;Q�U	9�KUwv1�02oRwvpat�-�T�ange�/;Uh`#C j80��WeldConGdMo���H�JK0�#7a�Dq (T����iJ\atk30�e���R�1�{�wm�]MON�_�0\��$�_��$Xg��p@��b��"At�<�%stop�/r�@����Zd��y8N4�Cir��ld P	r��XvF�ׁ��K
��1��cS7�O1��1\q�-\?8�at_ufrm.� #E�R�7xcArc A�bnr�l \it�ob9  �H552}�12{1 [prc���2 a�1AAgVM ��20 ��?J614��@�TUP mch �"#@545�PC�#B6��VCA�M awam�0C�RIMe_@UIF���#A28 0`vr�_@NRE�b.@R6s31�s�0SCH���DOCV l�isi
@DCSU�E�#A045pR51?EIOCe t���0542}�R�A9�6 pC
@ESEkT ��c
@J5K@���#@7K@;bM�ASK acry~v@PRXY cw1�wB7%��0OCO �Pht�B3�s;B2�  Q�B0�p paa#A@4�;A39�0�Fo�@H^SI�oLCHK�@59�@�OPLG ��;A0�3 ��PHCR �:�PCSP  G�W�R6 ��;A54���PDSW@_f��0MD;P "FO��@OP;P�PPR�O!ÏB7 mfo�rk�B0�UPCM�F	e�@4f507��U�@5-hg��!fR�ST-f69`cl�mPFRD@�SR�MCN	eH930ށeSNBA�USH�LB	eSM�`me�xte�B6�fPV�C-g2�`��~QTC�P�UTMIL	f7�895@ups�`P�AC�fPTX	eTWELNrd�R9Ef�8@w1 mpu�sh#@958Ef9{57	eUECKYu�UFR�fVCCM�	eVCOR	�k.�vS@IPLU�@I� ��_f�qXC ykZ�_@VVF �WEBP Y���aTP��t.�pR�626 T In�pCG�pnF��I=� ��6�PG�S�R3_q95 7�18 P�0738� f��1�@
  ���AC`6�A63 w794�B523�5�R65�1Sua5'53 ��A4�@gC�=@1qED064 /tamapF����O�6 sths.^_@LIO ��w^p~��5 - HefPOCMSC��ӂP���51@STYL <t�_@TOP ��P�R5{@Wave,��PRSR ���A8-01UOL�Ph� v@OPISY0��`� w.��0L�p}���S��t^pETS��fun�0SLM�TY0��B9 62�3�A�`E�5FVR�C�0_��NL t�j�wp001E��2�E��3)E��6 j���:@U0'@BDݐ5�MEݐ8 a֐��U�0�`6������5(��?@s@S���0�F�61�=�3 ���;��@69�U5�`*�faF�_�7 h��݁a�8Y�04^�!9��_�_PT�up���20w0��6u���71 ���@��8 �"���9u�us�0U�1a�w�㢸�{@Ʀ�@Ҧ3�3ݧ38`���`
��@�7 R.$ML��/�K ���9����40E[�1̀S�e�@]�2��Ea�A�NRSل� �33�4���拰��n�e���Roboz���net�����ደ��9���!拰j��\srvo���4�@h���x�����Srv���t ROB:PM'�e�4��5��G�n��r��b*ŋ�ite��ӿ�5�-���6拰35v��564x��7@Main��tatio����6@����������o����S��, '���t 拰\��\cc��? "TORC���`�����L��crV�CCR�����5'�xk965���� ��N���MО�6�����;���o_��w5�߆�0ch��y6���v!.j�k��iw2�߀
��x5�����2A.���n���3V��h�z��5���ui)f����c��_�3E@H��,�l�����T�1���T�2�(�Z�l�4z���?������/�l_i��}3Ѧ����0� |�{��  Y2�?�jog\dju�i���og��awWmfr� f��F� �ius�� Eq LibJ��6K񄐞S��/3�� (�bA,��2�7�_5'�\�<��� "MF�����d5a��n7y57eM��m K��߽Ҡm���g �����̞A�tw1������tw���#���6 'ink��0LR .ќ�6��J852���J�597�98��88�J�!�1^%N6���b�GN ��k\etl�@.�CO���O#|A` "ALNK
�>�%rd_�PB�� �"\wr*1O="�"lS ��P$d��0�88����PN A;RC��PRM�3��@B0��Nŋ��!8^�<���1SU P��$P��Ç�H���0��|pм3mpana/'p�ȣ0�1��H57X��85n������ �0K�BH@��<��1��bel������R��<D41��HDY�dhen��8<A���D���Cm���EN������D.��E��<�!� kemp��Dh¼3�m:re��2��pEf"sFMIG6�A00��37JR��|P�!�IGC (�P�.�E�%�чߑT� a;vs��IGE��Gџmigco`'�m�n&NA�ц�fa�vavtj�VTP�o/lfrm "S؆pGoYmsy�ASY�qo/lpdhV�PDyH�oYktpdl7�DL�o/lrf�`CRF�d�y�p8�3b:��s�`.vr3h1y�rLO5ccr��p �4c�§��q�@�����������R�RB�Sg�S����.�o���.��Z=fArbt\��`c.2  �w� _	b���! TertiB
ELS�P�2�U�g��YL (Co�mmyle s�eU�%)��bգ�s���'�ps01 "�PS��.#le\pscol���u.�6��ry�Pr: ���vׁ�Q�4syrs�r��-���ice Requ��g%���SRS�2K�9�P6k45.�9R S�"H|����(����vb�Ы/�,M�ۂfO� " ��s�O��sr������aP5A��+�m8���2813�P�49Z�89���A��{��Z�.���g�st�M�\����|�8
?�M�utl�v��'�&Q�N����q s�pdramj�!�peed.�pf%�Q���NN05���J67��2NĻ�� j�(��d� RH�-�	D��b ?"RMTX"��Ə~E�  ;�2 "S�0q�Q�D���slmt�o�ft� mi��SmL��H6Q64봷H62F�20�6c07B��P�38e��2 Hk�e�s�;�5�l�62K�79��7�95�79��60U9j�1F�1x�4��e5��2����H6���843[�2s�8215j��6�MT+�"�@��6����f�� "����S��\Af봆봖�0n��- Positi5o�l��esf �F�1N1h�ݻP(���ti��,봥�ǀ�ņn1Z�POS�s� �0� �h�873�r�riv�e Axes+�H�8��4di��(D�ual Dr�sHΕ�Ȅp��C�\B��j�.�kŔ*�ex�sj� De)�1��63����AM Indexjź��x�&�\ami:�s� �mi&�8�c�a�sC��nt Aongle+�CO;�p���봗#COM��Mom�������Ϋ�gou���! ̂�
fl���Envi� m���6k�d��820)����flx(�2� |�r��ionΓ{�ǅK�r772\ic�P�$	� �x0Z˱t;��2atzn������c�TJ�ync�Ins�p��R76��� �#���Xj�r#mSB����T�b5=mK�masyA`j�ܢ�nc\��MA�SIr�{��b�as��ulti-!A�`�6V��7v!� +��5k�NN�P ���se��!\��FGRLK��v�k��hdzՎF봅"fr�lk��&�m
ŊTr4���C��il/-&�e��r7��0Zo�nd ��:���� "ICRZp�%Q�g8�Piabic.]T�IAB0c���0o�e�I�0V�E �0��1 (�1�4���0濡�0�C�2\i�0t� IA˱�����"�@AiciAC@�0b��!�1�1��!�0omain�sDP�1�n C7`[��0e�DLPV�2�0��hpV��P M_@��̘ ��O]B�ưI:A��Єdp�CD�O�F"�0N>I�A�B���0_�Fd%4�e�o@nn Stan��A[�'"� MCNl�>�90�096:��s�5j��0�Q=���H��0���Q�2~Q(Re�m^PkAeSdard�I0��W2�NQ�0\t�prcmuǰCM�U�ku�1�TRP\r�c�0�q��jBRSUF1q73 �0uip��[��Ae�J61S 5�9Q�I�0taV"i Eq[A��Ζ�Rǅ�!2ȡjt`�Pcp���Esr��A�Qvb2 h�Q⦷ka�@xa�0 #�-���1 �a:��1� awmgenl��q�0ener��Woeld zQiboX^�0AWMG�U7{o _q(G>t�A�`%�b�;�d�60t[A3rt�1.y�R mshc�q@�3��n she�qqGR��1CMSC �U�A���RhjQ����p�0l�0rd$�1�8� p[a��u\qs�h� PSH��� �X  ������0   (�L r wKq�1/�Fe$�Q7�Ij��\;cl
A "J����0 H\j�Qcle���"E�S�Heӄu�ybU��`{A�ybm�dprm"�8�zal?i_varsS�돞��iconu���d�bg"��0Iz�ցrgpged"��1�&6��� Ԅm_�0�1x�i�Q҃m102؟��e_no��ȕw�rspq����wr�pirS�[q>��0gCas��Y��1��_s�ƅ�wr������ff<ӯE�inch30U�>��extwd�N��wrc����'�DՂrdS�Q��0"!�i�����aN�b �i����0�Ə(�/i@��RF�p
q���saj��ca��ntKCMAP ���O D�B�)��T�f�ap"Qj�AP�C��Z���0stmN(PSTM.Q{� ��apcevre*a�o��in
Au7a*a��is
�rbCIS�D G�QMete0/`�3�0T56��i�<�cQ��Q7�ar �>�,KQ�Y��(�\sl(�gr0S�14�e���q�	B..i�A������d��/�[a��>ֻ1���Q�d+Q�G 
�(5ф�M�Q�O K�џ� `+�2�`KQ�����B ��Kq��GT��sU�0���0S30le Ac	t�C�8R��Y
AQ�4.��1�㵏�I��-\J�ds��SU^� %����{A�#���s�!�j691.f�1S�ervoTorc�h9��6Jv�K� 91 (�K�A���Q�svt��VR��AsRC
�es4 F���Q4��MU�dq�v�z�vt/���5�+Q tFEv� ՛0"S`���0h for A�lumi��982Λ� 82������; ��	��d�L{���oo�q��l���L�ϊ��\srvt.vK�3e��0�0hP�AS`�� A��<^
�S016F�85�(�0�*�(!ez���hS�ATNQ���h`
�"P�QNG���	��2w�ADW����t��ҋ�М�wenmr�8sn�hanced M;ir�bmag ��b7R69�Q90�+�E.'KQ I>!��I�""\mjQr�MI)R�c;� � e$!.b�06b"%�tmbuswtcpy�Mod� / TCP��REˑX nvkAd�8���!K3CP>� \�$�P}m:1"MBUI2���i2d0� i�+�%���p�930�sPRO_FINET��OJ���J93+� �0 (�5��>鋁Y�3�P?pnio ":���x�1"P�q(@RIO��/ǖ$A��u�3)tj#96Od:��@gT�UHc67J�O��Q�`FSW䑡@���?K�67\fswpr��W+F�}�A\f_��ach޷	�A;be�r4���96�p_f�wd!6���f_r�ea/T[O 'Qneu4��_�Rr��sR��C�Qurn���%S�enא� $Ssw��t�_fswcol�#�n�AQ��Ak��cvvcuj�2�i�RCalib V~z!nc Utl4�OVCUT� ��1?��b(�a��VisF�u�cj���`k�vc�cU���c�tpfia�_z��`p6b�_8+�apset�3���c\z_�p{���k���uKA4���c��j9�88/�To��orYs1�!�p.�=8�?5 �p ^ol +!p��+��p\gf*��D�sT�c���V�Mas@��9�;� �|�����1� P�osij�����or�dt���v�
�02\���up޶�����r�_dc1$AB�As.��I[\N�bj An�e��b���򾿀��ۿ]���+�ޘ�� �_wQW�� k_Bc0y�t{G���F4�1�k�nifi3 sSpeY��94� a�1�UI n���v�>��k1��`�\frco���
�j9��1�Brake ch:ѡf�`0�{Q�5GJ��(�ck�rpȺ���˕51��b��BRCHUCD ����P�����5/�C����m�ulaneous��=���>55`�lo�H�SiɀS�TD u�LA�NG ��!�c�s��0C�T��\�cscsm���1ﳔsﳠ�=��C8ﳡ�N�dss' �Σ@c S�F�
������3�V68��F�,��sﳥ�s\��u�ߣ�ć��N�r69����gn�ost�eo� n������1�U�i -��9��C�ﳵ�7�z!�\�"DVMV����"r6�Đ�ﴃ! !��p��Uԧ� tr�D!ﳢ��2ﳡ�[�4� TcԦ���er�!��q>+�\pc3j��׸��Ƴ075.�os.Re���rN��� g��2c�6��ė�� �|����75\pt�TJC6���b���Ā���Bg�ė@I�>�S�i>��80��J979a�08� 1���(Iepi{�UL+�oﳔ#��a��f "NRU���¡�prsta�2�£��gutl.��RBT��OPTN�q0\?�r?V�@H nr?�ro�vq?l rb?r�DPN���!�r�rdfi���u𷁟�basi1c�ߡ�fc� ��J��A-�q��H�829V �$��9��@������Ph>�c "F2�
��29���j83���ce C�t�our� UPDT�3�5����Fo��on���aг�Ӵ�Q8�ho�ff���r� 35�fnV���r��\f�V�����\fcn��rg%3($��% ��r�A������6�%�D �E������g0@=��$���$n���/1!46%u��C/ T0\> ])A��av2tp�0ޖ�0v�0�2Av6`�0���0?U8�0 �1Br�0���0�4U0L�vpofs`1|��1|�3y0� mgp�s�0Nv�<un�Q�,x�0�4se�5ҌBT0�~�b cellf�1��el�0Cp���1©�R�1�f�B��51=9�1ll F�B�0@��p�0b�C�Bn�0/fncl��"RA���Z�0^V�Bfndrxu��AsIND"�1��>�A�1\fn��t��A^f�0t�B&PTPe�xjA�?�@�0%QTPc��1�v�1u�B&Ptqd~_�[ Q�2�V�G�j7��0- V-�500i/�010i 3D�0�[S ��15�`ab`�1�3DE��0N��<9\�calc@�_.27~�0vsfit3Ep �0�{a���07�u�0\`�`Tra�0B��KJ�a�MJ�`�b�e �1�bE��10Ov�0=j�`\que�1�?��3Arpo��8_�`8��1epush3��� ���0}s\�М�v��/�qkm�1ޕ\��swa�?�h�qaiynj|wkclb*O���?qvs
AJ\ud�sblt���ee�nn�g�|wigc�hk��uv�avu�A�s�� |���0  `�тv��3��_p��FA��GA"73�1c�ro����,�v�Apo ��0�8�a�jB���iR�qon E�rro9���.m�FQ�A757�Aж�1�� (iR�A���R�.]kZ�<d\mh/erhd�AH4P��<�}��\ire:AR���ree���/0�B�@���l��Z�h:Ahd��� ������j���cv�a���`�1SP APAS�A��SA�Sz�09 �q C�TAMڠQTABjڡP�AGz�13�Ҷ�Π(�`�Q�����p&u/M��pas\�aama�s+�=�
A`F��c��s��bia�B?����VS����VSIAС��D�q�����(�A��vA�C�  �6� ϼ���1 ? !   ��M� �Ó0(�8� ��\���>ұ(H� ��]ia\ia�`�a�`h���P�g�QoiZ�Ƴ|c�������  ����*SY�ST�EM�0A ����$ˢ�S  ��0����������ATSTKSI�Z������0����� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y������� 	-?Qcu� ������*��Ȳ��TART_�T SAG��$}D��IGNAL���SARTUP_CNfQ/a/s/�/�/p�/�/�/�(J�2!
�
 �/?? )?;?M?_?q?�?�?�?ܹ?�:99�$K���$FEAT�_DEMO C�����1@   �8MO  OMODOVO�OzO�O�O �O�O�O�O_
__I_ @_R__v_�_�_�_�_ �_�_oooEo<oNo {oro�o�o�o�o�o�o A8Jwn �������� �=�4�F�s�j�|��� ����̏֏����9� 0�B�o�f�x������� ȟҟ�����5�,�>� k�b�t�������įί ����1�(�:�g�^� p���������ʿ���  �-�$�6�c�Z�lϙ� �Ϣϼ���������)�  �2�_�V�hߕߌߞ� ����������%��.� [�R�d������ ������!��*�W�N� `��������������� ��&SJ\� ������� "OFX�|� �����/// K/B/T/�/x/�/�/�/ �/�/�/???G?>? P?}?t?�?�?�?�?�? �?OOOCO:OLOyO pO�O�O�O�O�O�O	_  __?_6_H_u_l_~_ �_�_�_�_�_o�_o ;o2oDoqohozo�o�o �o�o�o�o
7. @mdv���� ����3�*�<�i� `�r�����Ï��̏�� ���/�&�8�e�\�n� ��������ȟ����� +�"�4�a�X�j����� ����į����'�� 0�]�T�f��������� ������#��,�Y� P�b�|φϳϪϼ��� ������(�U�L�^� x߂߯ߦ߸������� ��$�Q�H�Z�t�~� ������������  �M�D�V�p�z����� ��������
I @Rlv���� ��E<N hr������ ///A/8/J/d/n/ �/�/�/�/�/�/?�/ ?=?4?F?`?j?�?�? �?�?�?�?O�?O9O 0OBO\OfO�O�O�O�O �O�O�O�O_5_,_>_ X_b_�_�_�_�_�_�_ �_�_o1o(o:oTo^o �o�o�o�o�o�o�o�o  -$6PZ�~ �������)�  �2�L�V���z����� ������%��.� H�R��v��������� ����!��*�D�N� {�r����������ޯ ���&�@�J�w�n� ���������ڿ�� �"�<�F�s�j�|ϩ� �ϲ���������� 8�B�o�f�xߥߜ߮� ���������4�>� k�b�t�������� �����0�:�g�^� p�������������	  ,6cZl� ������ (2_Vh��� ���/�
/$/./ [/R/d/�/�/�/�/�/ �/�/�/? ?*?W?N? `?�?�?�?�?�?�?�? �?OO&OSOJO\O�O �O�O�O�O�O�O�O�O _"_O_F_X_�_|_�_ �_�_�_�_�_�_oo KoBoTo�oxo�o�o�o �o�o�o�oG> P}t����� ����C�:�L�y� p����������܏� ��?�6�H�u�l�~� �������؟��� ;�2�D�q�h�z����� ��ݯԯ� �
�7�.� @�m�d�v�������ٿ|п��  � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r��������������� &8J\n� ������� "4FXj|�� �����//0/ B/T/f/x/�/�/�/�/ �/�/�/??,?>?P? b?t?�?�?�?�?�?�? �?OO(O:OLO^OpO �O�O�O�O�O�O�O _ _$_6_H_Z_l_~_�_ �_�_�_�_�_�_o o 2oDoVohozo�o�o�o �o�o�o�o
.@ Rdv����� ����*�<�N�`� r���������̏ޏ�� ��&�8�J�\�n��� ������ȟڟ���� "�4�F�X�j�|����� ��į֯�����0� B�T�f�x��������� ҿ�����,�>�P� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������� � �$�6�H�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
.@ Rdv����� ��*<N` r������� //&/8/J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�?�?�?�?�?�9  �8�1O(O:OLO ^OpO�O�O�O�O�O�O �O __$_6_H_Z_l_ ~_�_�_�_�_�_�_�_ o o2oDoVohozo�o �o�o�o�o�o�o
 .@Rdv��� ������*�<� N�`�r���������̏ ޏ����&�8�J�\� n���������ȟڟ� ���"�4�F�X�j�|� ������į֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*< N`r����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?�?�?�?�?�?O O0OBOTOfOxO�O�O �O�O�O�O�O__,_ >_P_b_t_�_�_�_�_ �_�_�_oo(o:oLo ^opo�o�o�o�o�o�o �o $6HZl ~������� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d�v������� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p������������� �� $6HZl ~�������  2DVhz� ������
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�?(�?�?A@�8O ,O>OPObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟ޟ���&�8�J� \�n���������ȯگ ����"�4�F�X�j� |�������Ŀֿ��� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�t߆ߘߪ� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: L^p����� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я�����*� <�N�`�r����������̿޿���$FE�AT_DEMOIoN  Ā2������INDE�X'�6���IL�ECOMP D����h��5��^�SETUPo2 Eh�r�?�  N ��[��_AP2BCK �1Fh�  �)�����%�����k���/����[��� �ߌߵ�D���h��� ��3���W�i��ߍ� ����R���v���� �A���e������*� ��N���������= O��s�&�� \��'�K� o��4��j ��#/�0/Y/�}/ /�/�/B/�/f/�/? �/1?�/U?g?�/�?? �?>?�?�?t?	O�?-O ?O�?cO�?�O�O(O�O LO�O�O�O_�O;_�O H_q_ _�_$_�_�_Z_ �_~_o%o�_Io�_mo oo�o2o�oVo�o�otwɫ�P�� 2��*.VRN�`*Qw�c}��e�8pPC���`F'R6:��~�"��{TF�F�X��uC����)�����f*.F�;ُ�a	�sǏ�x��*���STM J��S�^��pK����`�iPendant? Panel����H���p�ϟ���3���GIF=�g�r�S�p�"�����JPG����r�ׯ����;��zJSE�n��`�\���%
JavaSc�ript��ůCS����q�߿�� %�Cascadin�g Style ?Sheetsϐ`�
ARGNAME�.DTMϰlu�\�a�ρ��Ģ�N�	P�ANEL1����%�u���%ߜ�����2 ߀��n�+�=�����3�����߯���V���4"���v�3�E����Y�TPEINS�.XML��}�:\������Custo�m Toolba�r6��hPASS�WORD��nF�RS:\y�8� %�Passwor�d Config ���o����9�o] ����"�F�� |�5��k� ���T�x/ /�C/�g/y//�/ ,/�/P/b/�/�/?�/ ?Q?�/u??�?�?:? �?^?�?O�?)O�?MO �?�?�OO�O6O�O�O lO_�O%_7_�O[_�O _�_ _�_D_�_h_z_ o�_3o�_,oio�_�o o�o�oRo�ovo �oA�oe�o�* �N�����=� O��s������8�͏ \�񏀏��'���K�ڏ D������4�ɟ۟j� ����#�5�ğY��}� ����B�ׯf�Я� ��1���U�g������ ����P��t�	Ϙ��� ?�οc��\ϙ�(Ͻ� L����ς�ߦ�;�M� ��q� ߕ�$�6���Z� ��~���%��I���m� ���2�����h��� ��!�����W���{�
� t���@���d����� /��Se�����<N���$FI�LE_DGBCK� 1F��� ��� (� �)
SUMM?ARY.DG��OMD:!a� �Diag Su�mmarybo

CONSLOGW�:L��tCo�nsole lo�g�n	TPACCN�@/%(/e/p�TP Acco�untin/o
�FR6:IPKD?MP.ZIP�/��
�/�/q� Exc?eption�/�+�MMEMCHEC�K[/�Pq?�M�emory Da�tar?ra,])}]1HADOWg?�L?^?�?�3Sha�dow Chan�ges�?�-�?�)	FTP�MO��?QO|7�mme?nt TBDzOr�=t)ETHERNEToO�01��O�OtEthe�rnet �fi�gura?udADCSVRFnOTOfO�_�1%DP v�erify alyl�_�10"�?UDIFFw_]_o_o�0%�Xdif�fo�W01DPCHG�D1�_�_�_�o �o�o�S!�Gi2pofoxo �o4�oGD3�o�o�� #�Gv�UPDATES.��p��FRS:�\��uUpd�ates Lis�t��PSRBW�LD.CME����Y���PS_R?OBOWEL�Om ޏ�����8�J�ُ n�����!���ȟW�� {���"���F�՟j�|� ���/�į֯e����� ����T��x���� ��=�ҿa���ϗ�,� ��P�b���Ϫ�9� ����o�ߓ��:��� ^��ςߔ�#߸�G��� ��}���6���/�l� �ߐ�����U���y� � ���D���h�z�	� ��-���Q������� ��-R��v�� ;�_��*� N�G��7� �m/�&/8/�\/ ��/�/!/�/E/�/i/ �/?�/4?�/E?j?�/ �??�?�?S?�?w?O O�?BO�?fO�?_O�O +O�OOO�O�O�O_�O�>_P_�Ot__�_�_ � �$FILE_��PR�����P�����XMDONLY �1F�U�P 
 �;_o__6o�_Co lo5_�oo�o�oUo�o yo �oD�ohz 	�-�Q��� ��@�R��v���� ��;�Џ_�����*� ��N�ݏ[������7� ̟ޟm����&�8�ǟ \�럀���!���E�گ�i����ZVISB�CK�X�Q�S*.�VD�a�ϠFR�:\0�ION\DOATA\L��Ϡ�Vision VD file�� ��տ������/Ͼ� @�e�����ϭϿ�N� ��r�ߖϨ�=���a� s�.ߗ�&߻�J����� ����9�K���o��� ��"�4���X������ #���G���X�}���� 0�����f����������U�ZMR2_G�RP 1G�[�C4  B�> �	 �Q��� E?�� E�@����`
� OHcGP{�K���/Jk��?� �`� :G:�<9�{��H�A� � dvBH�C�{�N�B�ƈ��`�� z  �D���>��	@7UUU�UU�`�/���#@=u�dѽ��H=���=�~�=��yC,���;��.;!�9����:�b:�l?��/ /�/�/��E�  F,D .�!D�`�#�u�-ދ�E�� �!D+�2C�dR_C�FG H�[T ��/O?a?s?�N�O �X��
F0�1 �0 ��  �0��PRM�_CHKTYP  �P�> �P�P�P���1OM�0_MI9N�0<���0�P�X�PSSB%3I.�U�P�#O�:CCOUO�UTP_?DEF_OW�P:��YpAIRCOM��0{O�$GENO�VRD_DO�6��R�LTHR�6 dz�Ed�D_ENB�O{ �@RAVCx9JGC� ��[OF_�/j_�x_�_7��P�QOU{ P���B�8�(�_�_�_o^o  C�f`\Voh�X�oYm%~oBȽ��b�	�Y\OPSMT�SQY� @ed�$�HOSTC%21R�9��G�  5M:}k;8  27.0�p=1t  ek� ����z��1�C��U�x|�	�	ano?nymous|������Ώ��7:� �� ��ik�P��t����� ����������9� ӟ��^�p��������� ��+�-��a�6�H� Z�l�~�͟����ƿؿ ��K��2�D�V�h� ��ɯۯ����#��� 
��.�@ߏ�d�v߈� �߬��������� *�yϋϝϯϱ�{��� ���������Q�&�8� J�\�n������߶��� ����;�M�_�q�F�� ��|������ �0S����x �����K!3/ Gi/P/b/t/�/� �/�/�/�/�//Se :?L?^?p?�?��� �?	?�?=/O$O6OHO �/lO~O�O�O�O�?YO '?�O_ _2_D_�bq�ENT 1S�[� P!�O�_�R  w_�_�_�_�_�_�_ o �_,ooUozo=o�oao �o�o�o�o
�o�o@ d'�K�o� ����*��N�� G���s���k�̏���� ����׏%�J��n�1� ��U���y�ڟ������ӟ4���X��QUICC0e�A�S����w�1�������w�2����T�!ROUTERU�1�C���!PCJOG�����!192.�168.0.10�~�s�CAMPRT,��ѿ!�1���RTn� �2ϓ�YTNAME !fZ?!ROBOϛ��S_CFG 1R�fY ��Auto-sta�rted�4FTP�?,��?�OW��? {ߍߟ߱���hO���� ��@�.���e�w�� ���6��)���=� _��F�X�j�|�K�� �����������0 BTfx�?�?�?� ���3�,> bt����O� �//(/:/��� �/��/��/�/�/ ? ��/6?H?Z?l?�/�? #?�?�?�?�?�?K/]/ o/O�?hO�/�O�O�O �O�O�?�O
__._QO R_�Ov_�_�_�_�_O O1OCOE_*oyONo`o ro�o�oe_�o�o�o�o o�o�o8J\n� �_�_�_o�;o� "�4�F�X�'|����� ��ď�i�����0� B�����ɏ��� ҟ������>�P� b�t�����+���ί������T_ERR� T���"�PDUSIZ  ���^ɐ�9�>R�W�RD ?�Ō���  guest��������ȿ�ڿ쿣�SCD_GROUP 2U�̫ ����1��!x��2�ǒ  ,C��	$SVMTR_�ID 2�Ti��$GRP_2�$�AXIS_NUM� Y�z�f�NF���SV_PARA�Miɑ� ,$�MOT_S��TT�P_AUTH 1�V1� <!i?Pendan����Jũ���!KAREL:*��݇KC3�C�U�+��VISION SCET��ߊ���!�� ����(������e��<�N��r����CT_RL W1������
��FFF�9E3�FR�S:DEFAUL�T�FANU�C Web Se/rver�
��z� ���������������� �WR_CONF�IG X!��m��"�IDL_CPU_PC0����BȊ�K  BH1MIN<)�OGNh�O+�`���7��3 NP��IM_D�O��TPMO_DNTOL� �_PRTY�K�OLNK 1Y1���#5GYk|}�MASTE� ����	OSLAV�E Z1����O�_CFG��UO�����CYCLE���*�_ASG s1[l�
  ]/o/�/�/�/�/�/�/ �/�/?#?5?G?�0"ď�`�5�_��IP�CH/���RTR�Y_CN0���SCRN_UPD_���9� ����\1�&�O&��$J�23_DSP_E�NB�01�%�@OB�PROC%C��J�OG�1]1��8��d8�?�R;�OR??U�S��LQ�O�O_#_�OG_Y_�k_}_��'ҟ_[CP�OSREEO�KA/NJI_�K��S$1��3^���U�_�UCL_L[ m2�?��PEYLOGGI�N�&��}A9���$LANGUA�GE m��2*� �a"�LG�2�¬������x&аҘP���Q ���'0ꩨ����MC�:\RSCH\0�0\�}`N_DISP `1�����8�O�O �LOC�B�Dzj�A�cOGBOOK a;+�~@����q�q�pXCy�����*�b=�0�O���	�u��y��Fu����!ua@B�UFF 1b ��2��ڏ�r���� ���$�Q�H�Z���~� ������Ɵ������ �M�D�V�����DC�S d�} =���L�����!������!���IO 1e�;+ 
OZ���� Z�j�|�������Ŀֿ �����2�B�T�f� zϊϜϮ����������
�5�Ez TM  2{d�_c�u߇ߙ� �߽���������)� ;�M�_�q�����8��qw8�SEV�02}]4�TYP@�R�`3�E�W���QRS? �Ko���2FL 1fC��0�˯������`%7h�TP_`�@�"�k}NGN�AM%D�e���UP�S*pGI�5a�5��_LOADB@G� %2z%
OUVREPINC�0���MAXUAL�RMm7�{8�_PR�4�0�sM�C-pg;)[�q�sx�Pc@P 2hV� ��	"��
�0���t��� �� /ɨ/O/:/s/ V/h/�/�/�/�/�/? �/'??K?.?@?�?l? �?�?�?�?�?�?�?#O OOYODO}OhO�O�O �O�O�O�O�O�O1__ U_@_y_�_n_�_�_�_ �_�_	o�_-ooQoco Fo�oro�o�o�o�o�o �o);_J� fx��������7�"�[�D_L?DXDISA� B��3�MEMO_APދ E ?��
 �c���ɏۏ�����#�5�ISCw 1i�� �M� ���b����L�՟�����J�C_MSTR� j���SCD 1k����g�� ��v�����ӯ��Я	� ��-��Q�<�u�`��� ����Ͽ���޿�� ;�&�8�q�\ϕπϹ� �����������7�"� [�F��jߣߎߠ��� ������!��E�0�U� {�f���������� ����A�,�e�P��� t��������������+O:s	�MK?CFG l'�n~�LTARM_�m���q����,METPUl9d��/�ND�CMNTd�% � n'�c���{�%POSCFz1<PRPM0��STOL 1o�'� 4@C�<#�
�n�/'� //1/s/U/g/�/�/ �/�/�/�/?�/	?K?�-???�?k1%SIN�G_CHK  ��t�ODAQ�p�=���5DEV �	'�	MC:>�<HSIZE��C��Ȼ5TASK �%'�%$1234?56789 \OnE��7TRIG 1q`��%H��OA��O�O�O)�>FYP)A�E�4��3EM_INF� 1r� �`)AT&�FV0E0�Og])�OQE0V1&A�3&B1&D2&�S0&C1S0=>V])ATZg_�_�TH�_�_vQ�Oo�XAo?o�_coJo�o�o M_�oq_�_�_�_ �_<so`r%o�Q �����o�o&��o �o�on�y3���ȏ �������"�	�F�X� �|�/�A�S�e�֟�� ��1��0��T��x� ��q���a�s�䯗��� ��,�>��b�����A� K���w��ǿ��ɯ :�����#���G��� ����ϡ����#�H��/�l��?NITOR�LG ?K   �	EXEC1Tj��2��3��4��Q5��@��7��8��9j��6���� ������������ ����������U2!�2-�29�2E�U2Q�2]�2i�2u�U2��2��3!�3-��3�һ1R_GRP�_SV 1s<[� (s1�$���<?�lk��ʏ$�c�ڌ�=FA_D�,N�P�L_NAME �!S���!D�efault P�ersonali�ty (from� FD) �RR�23� 1t)4��x)4�����0@ dp*< N`r����� ��&8J\n�82���������
//./@/�2< �j/|/�/�/�/�/�/��/�/??0?B? �  �\  ��  ��`���  A�  B�m0Tm0��0
Y0��]0����  ���i0h0Bm0pm0ȷ  C�0C�0P� D�  D����2E@�2�2z �0�1�0�1�2�0�9�2��0�6�4EK  E?+� E��6�2`�0�2 A DJZ��3 A@DI�2�5�4�9�:�1;�7�:�5�@�5�O��;�O�3�1�1E�1�~�0�` E���G.�4E���C�@Q��A] Y$UP�5#V� �DQL]hT�FQ8@�B  UA U�T�R YU Q|UU�@�Y�Q�]�Q �Y�@B�YAP�1�R 4oBg�UXo�S�1Q`o ng�Q�o�o�o�W�o�o �o 2DV`tU0�D�ΥE���orT1T1O�  l0��{q�d�s�t� �y���tpI<Z*����y����`q��0 b�-T� @�5?h0p��T�?q�p�q�@u���5o���;�	�l��	  ����p�XJ�����X � � ��, �ނO�K���K�zK����K@0>KH�K$�������趂�5��N�?��=P�@'�6\�����"��Iڿ��
��}v��?���X�������0�
=�ô�0�0���  �>ڃ���#�^���l�Y"�0���q����͔��'���h����i�� � �T��  ��`��v��	'�� � ��I� �  �-`��:�È��È�=���إ$�@���Z����Z�!�t'�5�o�N��j�O  '��O�@���?��@�t˅@��@����X���B&d0Cf�0��B�1��}q��C%
���. � W ��^�/�AB-`���$Ń��� ��A�q��1ș_φ�o�p�πϹ� �
�`�����n� �x��ݱ�� ؀��:�m�����?�f�f��0��� ���d�v�%��ߛ�?KY����|��(q���P�����ȃȄ2��?33�������;���;���;��D�;�$;?�< J]���G>Oހ�Z���=�?offf?��?&z�ޡ�A���@�,��j��u၄�� p���n���^約O�$� �H�3�l�W���{���`������+���F�p ��&��J��k��=,�ɘD�@����0�  F���� ��5 YDV �z�ƚG���/ a'/�N/�r/�/�/4�/G�A�0����O�tp��B�0h/?d/%? ?I?4?���pA�0t2 -`|1�?�u�?\?�2;�<��Ŝ?���?�?hOO*�į��W*O�C��@�` Ca'O*�4��0�1�A���ܨ���C>�CR BA��Aˉ7࢙���"���z���q��=��\)xO� ʊ=��=qA�B)�{���O� ��(��g�/P�q�Bp���{���8R��K����J?&DK���	HwW�H�'���!��LA�L��9K��4HŀHH� h_�zP��Lm��J�sdHK� ?H-�A��_wO �_�_o�_%ooIo4o moXojo�o�o�o�o�o �o�oE0iT �x������ �/��S�>�w�b��� ����я�������� =�(�:�s�^������� ��ߟʟ�� �9�$� ]�H���l�������ۯ8Ư���G�$��� C���4�F@��8��u�8�V����������Ͽп�����?��F( Q�`���G� ���x�8E��Y��>x�	3Z�q_�Ϧϴª�����ϰ�fC3�g����̅��?�3�Ȭ�ـX�F�|�jߠߎ��5P��P������N�`����.���P�0b����7���
C@�C@5����
� @�.�d�������������������������&  ?JK  �@^���v�����2 wD�J�E����0��B}1q1}0C)�f@�AC@@�?CB�J�J�m��C�����z���3��E�(��F���
/�/**@9$���4�C@C@���4�;
 */�/�/�/�/�/ �/�/??/?A?S?e?�w?�J�2��������$MSKCFMAP  D� �g!c!�>�3ONREwL  s��1��а2EXCFEN�B�7
�3�5AFN�CODJOGOV�LIM�7d@Bd��2KEY�7eE��2RUNULeE��2SFSPDTY���FE�3SIGN|�?DT1MOTWO�A�2_CE_G�RP 1zD�3\,�;_$�__q_� [_�_S_�_w_�_�_�_ o�_oPooto�o=o �oao�o�o�o�o�o :�o^pW�K�������1QZ_�EDIT�D�7�3T�COM_CFG 1{�=r&I�[�m�}
)�_ARC_B���DIUAP_C�PL��(DNOCH�ECK ?�; �������
� �.�@�R�d�v����������П����;NO_WAIT_L�Gl�	PNT1�|�;zi+F�_ERRQs2}�9�ф �����ï���3���^ńT_MOt�~{�x �>�D��8�?\_�I��b 6�m�PARAM:u��;�f&4����w� =� 3�45678901 '�9�K�"�j�|�Xψπ���Ϡ��������w��,�>�ѿb�ƃUM_RSPACE�?�R�o��ߥ��$OD�RDSP���F$HO�FFSET_CAqR�����DIS�����PEN_FIL�E��Ao����PT?ION_IOvO�A�;�M_PRG %��%$*t���WORK �W'C ���6���2���S���	� �a���6�C����RG_DSBL'  DCj,@����RIENTTO��0���2 ��UT_SIM_DC���2�2��V��LCT �P�����>��_PEXE���GRAT��\F$E��>��UP ���x E �/A'es	��$��2St)4��x)4����@ dRߺ�� �&8J\n ��������/"/a�2�R/d/v/ �/�/�/�/�/�/�/��<A/?0?B?T?f?x? �?�?�?�?�?�?�?������)P�  ��  �p�A� g B!@�B�Y�@H@�  ���@p�B!@p�!@�d�c���P �D�  D��NbBE@jB_Bzd� `A`@{A{Bx@�I{Bd@��F|DEK  E+� E��F�Bx@0kB�A�D�JZ�fC�A �D�I�B�ElD�I�JlA;eGJ�E<P�Ec_}KPs_aC[A{AEhA�m@?�` E���WxDE���S��@�Q�Q@�]�Y�U�P�E�V��T �Q md�V�Q�@�R�U �A�U@dcb�Y�U�Q0e�U˵@�ida�mda\i <P�B�i�A�P[A�b�o �g�e�chA�Q"w da4Bp�gx�� ����
����"�A @E�W���P�s� ��j�����(�(��� �O 1y(�Ho(�&��`�o0��C @�Eo�o��?|��C@�E��.�  ;��	lo�	�� ����p�X̰��q���X � � ��, �����H����H��H�P�uHV�2H�H_3��<���&��B�!@	�C����@�γ�4@L@�/
=�g��`@D��(�:�L�)�Aß�w½��ªV y�H@����p�ˣQ��֡�hD��D��  �  �������Q�6�%�	�'� � T��I� �  y��`R�=���x���(�@�������ʿ;��$�߯�r'�Np�"�  'F��:ą�Ca�B@CfBd�B�Au�G�Y� ��  ��C%�  ���^
��/V�B�`��p���;� ������wA ���^�'�M�8�qߨ��
�`��U�n� �x������ L����:O���Q��?�ffǏ���� z߶�%�ㅡ8��E�.S�?Y����4�|�	(����P���ő�������?333Q�����;��;����;�D�;��$;�< J!l�����6�޳8����?fff?��?y&2�A�D�@�,P�Q���-� 9�T�(���&����l� ����� ��$H 3l~i���� ��s������V���Dڹ@�U�@�  Fg�D��� ���/�/G/2/ k/�����-]/�/�/ =?y/*?<?N?`?��AL@��j��	�d�B8@ ?�??�?�?O�?B�'�A�*D�`4A ;O�0�?bO����S�}�?�؏O�O�O�O�Q��g��W�OC�>�P�` Ca�O�*�D��@�ALQ@I�	�b���C>�CR BA��Aˉ7��Q���"���z���q��=��\)0_�0ʊ=��=qA��B)�{�녨_�0��(��g��P�q�Bp���{���8R�MK����J?&DK���	HwW�H�'���1�MLA�L��9K��4HŀHH�  o�2`��Lm��J�sdHK� ?H-�A�Jo/_ �o�o�o�o�o�o�o %"[Fj� ������!�� E�0�i�T���x���Ï ���ҏ���/��?� e�P���t�����џ�� �����+��O�:�s� ^�������ͯ���ܯ � �9�$�]�H�Z���8~����KG�$��ſ� C�����@��8?�-��V��7�>�w�b���ψ�r������ϲV(xA�`����ϸ���0��ų�Y«N0߲S3Z�q_L�^�lҪ�x���߰�fC3�g��߶܅��?�3�Ȭ���ـ���4�"�X�F�EP��P��!�/���`�������`���0�S�>�V�7`�r�
{�{5��V����� ��������/I ��JXj�t��̪�����  ?JK  ���@.dR�r�2 wD��E���0�VB5A)A5@C)�P��A��@9O�X/"/2,C����2/�[/i*�CN�E�(�VF�i/�/�/�/R�*@�$�XxD�����O�|D�K
 �/E?W?i?{?�?�? �?�?�?�?�?OO/O�ZB��\������$PARAM�_MENU ?��� � DEFP�ULSE;K	W�AITTMOUTޓKRCV�O �SHELL_W�RK.$CUR_oSTYL�@�L�OPT��OPTB��O�BC�OR_DECSN�@{�N\H_Z_ l_�_�_�_�_�_�_�_��_%o o2oDomohAS�SREL_ID � +�x�@}dUSE�_PROG %�wJ%io�o}cCCR�@+�C�g_HO�ST !wJ!�d#�jT���o?s�qAs{�k_TI�ME�B�f�eh@GDEBUG�`wK}c�GINP_FLM1S�~�xTR��wWPGA � �|N���CH��xTYPEtL� hobo�� ����Ώ��	���(� Q�L�^�p��������� �ܟ� �)�$�6�H� q�l�~�������Ưد����� �I��uWO�RD ?	&�	�RS��PNeS��D��JOQ��TEbpF�TR�ACECTL 1���A ���� �e���� ߾��DT Q����ӰD ȿ 
 �����Ď`!�����	�

����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~�����z�����# 0)0 -?���������� ew������ �+=Oas �������� ;_/q/�/�/�/�/�/ �/�/??%?7?I?[? m??�?�?�?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�_ �_�_�_�_�_oo+o =oOoaoso�o�o�o�o �o�o�o'9K ]o������ ���#�5�G�Y�k� }���[/����͏ߏ� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� ���������!� 3�E�W�i�{������� ��������/A Sew����� ��+=Oa s������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?�?�?�?�?OO1O COUOgOyO�O�O�O�O��O�O�O	_Q�$P�GTRACELE�N  Q  ���P��'V_UP �����VQ^PBQ�WP'Q_CFG �VU@SQgQ���T9P�_�\kRD�EFSPD ��v\Q9P�'PI�NnPTRL ��v]P8�U�QPE�_CONFIrP�>VU�VQ�T��Y'PLIDoS��v]�QEaGRP 1��g���Q�C%  �ᙚ�QA�=qGY�� GcX Fg@� A�  D	��T	�Pd�T�i�i�5a5`� 	 p�_�R�[�o ´s�o�kBp>q�T>x�rH9B�!����~� �<T��<]/ ����U�@�y�d� �������я��⏠`z�%�P
�M��� ]���n�����˟��� ڟ����I�4�m�X������!Q
V7�.10beta1��V @�p��@z=q@��R|�aʡC  C5P{B|ܣDf@ ��C�`� D��� D� C��`�`B�䠃`C/�`p�R�r�`1��C�U�$�BdKNOW_M  �U~VBd�SV �mi�-e:�ſ׿� z����
�CσR�mAc�Mfc���8Plڢ	<�Rܡ  �b�� ^����S��ˠ`����I�iRLMRfc�Jy�T�z��QCz�`���u8�J�6mSTfa�1 1�V[
 0a-e��$բ�  �� �߽߫�������4�� )�;�M��q����� ���������T�h��2s���Q�<��a�3r�������l�A4��������l�5"4Fl�6_q��l�7����l��8�!3l�MA�D3V ^Vh�PARNUM  V[q2πj�SCH� ^U
�� )@S%UPD���e\/�_CMP_o�3PWP�P'WjS_ER/_CHK�%|X�&�/�+RS�}�Ba_#MO��/�%_�/\e�_RES_GrВv� ��nr?e?�?�? �?�?�?�?�?OO8O�+O\OOO�_44q�>< N?�O35��O�O�O53  �O�O _53^ _:_ ?_53� Z_y_~_53�  �_�_�_53K�_�_�_52V 1�v�$1���@c���"THR_INR0"!W�z(5dkfMASSxo� Z�gMNwo�cM�ON_QUEUE� �v�	6#0/�*�TNy U�!N�f�+��`END�a?yEcXE(u> BE'p|	�cOPTIOw�&;�`PROGRAoM %�j%�`�6o��bTASK_�I�o~OCFG ���o���DA�TArÖ�@0�2��t��������� g������(�ӏL��^�p���5�INFO
r×Q���d=�ڟ� ���"�4�F�X�j�|� ������į֯������0�B������Q� �lI�� DIT �����5�WER�FLIx^ci�RGA�DJ ���AЋ  ��?#0�d�R�G�a��y���?���a�<@���ɖ%ah�ϸ���[2����`\hF�]b2�2�A(dɻt$��*��/�� **:��#0��d��v���������W�Ab5�Ac	� �-�?߬�c�u߇ߙ� �߽�����N�I��)� ;��_�q������ ��������%�7�I� [�m������������ ����!�EWi {�����/� ��Sew� ������// +/U/O/a/s/�/�/�/ �/�/�/�/??'?9?K?]?�? 	 ��?�? O�7��9O��OfOO��O����PREF S�%�OpOp
۵?IORITY�g�}�߱MPDSP�q�Ϳ�GU�g��ڶOG��_TGʰ�r�j*R�TOE�`1���� (!AFs`E��`s_~W!tc�p~_�]!ud��_�^!icmX�_8o+QXYà��;�Oq)� ��2oDoOp�,omoPe\o �o�o�o�o�o�o�o �o;M4qX��	*)Sâ�MU������?&Ƽ7��/���K�V��~ȁƺ��AG�,  � �@w�������͏�E�t­C��O�Cղ߱PO�RT_NUMS����߱_CARTREP�@�����SKSTAW �J�SAVE ���	2600H738҈O�Or�*`������LÉ7�����7Z�URGE�_ENBʹ��aW�F(�DOV{�EVW�lPI�ձ)�WRUP�_DELAY ����=�R_HOT %�ֲ=�ɯZ��R_NORMALਨ򲸯�ܧSEM�I��Q���QSK�IPȓ��� x }O��yO��̿޿���= ϱ���4�F�X��|� jψϲ����Ϝ����� �0�B��R�T�fߜ� ���߆��������,� >��b�P����p������(�2��?$RBTIF7_�A�RCVTM[BT]�E�DCRm��t�� Э�E���A ELlC��e�@���8��o����O��ŀ��Aê|�r�5�9��]�顿��� ;���;���;��D�;�$;�?< Jl��Se ����� ����	-?�Q�GRDIO_T?YPE  ϝG�]EFPOS1 {1���
 x?� �Z@�</�^�� /v/a/�/5/�/Y/�/ }/�/?�/<?�/`?�/ �??1?C?}?�?�?O �?&O�?JO�?GO�OO �O?O�OcO�O�O�O�O �OF_1_j__�_)_�_ M_�_�_�_o�_0o�_xTo��2 1����oJo�oFo�ojo�3 1��o�o�o��o`K�S4 1�+=w��|��S5 1��������u���,�S6 1�C�U�g�����
�C���S7 1�؏���6�����؟>V�S8 1�m�����˟I�4�m��SM�ASK 1�z p�������XNOw⩦����MOT�EL�۫��_CFG ��b����PL_RANG��O�Q�OWER 崷��#�SM_�DRYPRG �%�%�����TA�RT �|�ʺU?ME_PRO�����&��_EXEC_�ENB  ĄW�GSPD��A�IȜ��X�TDBd�v�R�M��v�MT_��T�w��E�OBOT�_ISOLCخ�F�2�b���NAM/E ��É�OB_ORD_N_UM ?|���H738 �~  ����r����y� ��2�Dr�h�z�}�r� ����r�����
r��x�+��PC_TIM�Eg�S�xE�S23�20�1�����L�TEACH PENDANi�,����7���PM�aintenance Cons���$�"��TKCL/Cٰp������o� No Use��N��9ߎ��NPO��^����Y���CH_�L�����	�=��MAVAIL�SѸ�K�����SPACE1 2�� �K�����2�ļ�K�L�b���8�?����� IjAz������ ���':�_ pW������ �S'/:/�_ p/W/�/�����/ /#/?6?�/K?l?S? �?�/�/�/�/�/�?? 1?3?�?GOhO?OQO�? �?�?�?�?�OO-O_ }OC_d_v_]_�O�O�O �O�O�__)_o<o�_ a_roYo�o�_�_�_�_ �oo%o8�oMn U��o�o�o�o�o�o �z�I�j�A�� ��������/� !��E�f�x�O�a���2������͏ߏ�� �%�4�U��j���r�����3��Ɵ؟��� �� �B�Q�r�5�����������4ѯ���� �ǿ=�_�nϏ�RϤ��Ϭ��ϥ�5� �� $�6���Z�|ϋ߬�o� �������ߥ�6�� /�A�S��wߙߨ���@�����������7(� :�L�^�p��������������1��8 E�W�i�{���;���� ��9 N���G �e tE�
� �  e���// %/7/g�V-�c�/+�/�d� ���/ ??&?8?J?\?R/d/ v.g:�?�;�?�/�/^? O*O<ONO`OrOh?z? �?�?�?�O�O�?�?~O 8_J_\_n_�_�_�O�Op�O�O�O�_ `F @� +e�/9o_Ywa�Uo�o�o�_ zj{o�o�o�o I[%/As�w ����!�?��'� i�{�E�O�a���Տ���\
Yo*���_MO�DE  e@�S �e��_�ZA�Uo~�П��	��� �CWORK_{ADP�
xȡ/R  er g���Q�_INTVA�LP���[�R_O�PTION�� �[��V_DAT�A_GRP 2�,�XpDPP�� ����C�1�g�U� ��y���������ӿ	� ��-��Q�?�u�cυ� �ϙ��Ͻ������� '�)�;�q�_ߕ߃߹� ����������7�%� [�I��m������ ������!��E�3�U� {�i������������� ����A/eS� w�����W���$SAF_DO_PULS;�X��A�Z�1!CAN_T�IMO�!U��BR� �(�C�(��f0/������Ē����S  �����//��7/I/[/m//�/���C,"2�$��d�(�!�!�&�@�\
??.?*��)�/� ߠC4�_ 3b  Tf�W?�?��?�?�9T D���?�? OO$O6OHO ZOlO~O�O�O�O�O�O��O�O_�����%_X_j_'Y+a���Q;�o*����p(]
�t� G�Di�� -��,"���Q��y�_ o o2oDoVohozo�o �o�o�o�o�o�o
 .@Rdv��� ������*�<� N�`�r���������̏-��T?����+�=� O�a�s���ԏ�%��ß ՟�����/�A�S�X���-�0R2�S�U�] ����ȯگ����"� 4�F�X�j�|������� Ŀֿ�����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t�ߏ�ߪ߼������� ��(�:寧^�p�� ����������Y��� ��,".�@�R�d�v��� ������������	 '9K]o��� �����#5 GYk}��������X�$_�3/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q?�c?q:0/z?�?�6������?�=	�12345678��R !B�P

�8. �PO)O;O MO_OqO�O�O�O�A// �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_m�O$o6oHoZolo ~o�o�o�o�o�o�o�o� 2DoBH U}������ ���1�C�U�g�y�x����k;�j�� ӏ���	��-�?�Q� c�u���������ϟ��
iD���%�7�I� [�m��������ǯٯ ����!�3�E�oi� {�������ÿտ��� ��/�A�S�e�wω� ��Z����������� +�=�O�a�s߅ߗߩ� �������߰��'�9� K�]�o������� �������#�5�G�$@d�v�[��������)"Cz  A}�*   �(�2�4A��A!�
�0Ě22b�I[m,���0/���8���!3 EWi{���� ���////�S/ e/w/�/�/�/�/�/�/ �/??+?=?O?a?s?��?�?�?�?�$SC�R_GRP 1��(ӈ�(ӑ �@tw �
 ��1 	 �3 AB	D�� "M�7GJO8OqO���� nBD�` D��C�GnK��R-2000�iB/165F �567890. ��DX. R2D7� �@B#
123�4�EAFnA� CV�1B&�3�1��nAJBATY	�ER�_�_�_�_�_�\��H��0�TG�2&o5O6o\ono=FM/
Io�oEo�o����o��h,P�T~K� I�AB����B�ffBǿ33B�  +v��5wAA��G  @�
 _uA@�@o  ?��wrH-p�Jz�AF@ F�`x�r�=GC�  � �� ��D�/�h�S� ��w�7q_q�r������ʏ܄B���0�� T�?�x�c�u�����ҟ �������*��CZOH�m���  j���
�q@�r�O��=G��4߯-p���W\NCa�5�B$A�G�1Z�$�o�e �Y�
A {�����º��׸����Ŀ P�(�!�'�9�K��1EL_�DEFAULT � XT���
 _�MIPO�WERFL  t��w���WFD �n� w�^�RVE�NT 1����`u���L!D?UM_EIPM�����j!AF_I�NEk��B$!FIT��>��b�!"o·� �Q߮�!�RPC_MAINįߖ�������VI�S�ߕ	���F�!�TP9�PU=���d�5��!
PMON?_PROXY����Ae����Y����f���*�!RDM_S�RV+���g�v�!#R!T����he���K!
��M����i���!RLSYN�C5	8��Z!�ROS�ρ�4�I�!
CE[�MOTCOM���k���!	�CONS���l�>u�b9� /A��w��� �/�@///+/�/�O/a/Q�RVICE�_KL ?%��� (%SVCPGRG1�/:�%2?D?� 3+?0?� 4S?DX?� 5{?�?� 6�?�?� 7�?�?� TO<9O K�$��HO �!�/pO�!?�O�!E? �O�!m?�O�!�?_�! �?8_�!�?`_�!O�_ �!5O�_1^O�_1�O  o1�O(o1�OPo1 �Oxo1&_�o1N_�o 1v_�o1�_1�_ @B1�_�/�"� �/�  ��1����� @�+�d�O��������� ���͏��*��<� `�K���o�����̟�� ���&��J�5�n� Y���}���ȯ���ׯ ���4��X�j�U��� y�����ֿ�������0��Tϖz_DEV� ���M{C:\� 
�n�OUT`�h��j�?REC 1ŭuh��� �� 	 A\�������3��lu:��c�n�
 ��Tpvj6 s~S��  �����  �  �Пл�u��X�rU 1��h�=h����V�� ����h�+h���2������� ��'�M�;�q�_��� �����������#� I�7�m�O�a������� ������!E3 UWi����� ��A/Qw Y������� /+//O/=/s/a/�/ �/�/�/�/�/�/�/'? ?K?9?o?�?c?�?�? �?�?�?�?�?#O��� O)OOQO�OuO�O�O �O�O�O_�O)__9_ ;_M_�_e_�_�_�_�_ �_o�_%o7oo[oIo omo�o�o�o�o�o�o �o3!WE{� o������� /�A�#�e�S���w��� �����ŏ����=� +�a�O�����y����� ߟ͟���9��I� K�]���������ۯ��޽�V 1��� (�ӯ&���TOP10w 1���
 ���,�v�����@�YP�E��l�HELL_?CFG �{�h�=	�  ��B�RSR��/� h�Sό�wϰϛ��Ͽ� ��
���.��R�=�v߬�ߚ������%@�����ߨ������1������װ��2h�d����϶HKw 1�ݻ 
� ������������� ��+�=�f�a�s������������h�϶OM�M �ݿβFTOV_ENB����ƺOW_REG�_UI=ͲIMW�AIT:��mO�UT^�o	TI�M^���VA�L~p_UNIT�9�ƹLCW TR�Y^Ƶ��MO�N_ALIAS k?e	�he� Vhz����R� ��/�%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?�/i?{? �?�?J?�?�?�?�?O �?/OAOSOeOwO"O�O �O�O�O�O�O__+_ =_O_�Os_�_�_�_T_ �_�_�_oo�_9oKo ]ooo�o,o�o�o�o�o �o�o#5G�oX }���^��� ���C�U�g�y��� 6�����ӏ������ -�?�Q���u������� ��h�����)�ԟ M�_�q�����@���˯ ݯﯚ� �%�7�I�[� ��������ǿr�� ���!�3�޿W�i�{� �ϟ�J��������Ϥ� �/�A�S�e�߉ߛ� �߿���|�����+� =���a�s���B�� ���������'�9�K� ]�o������������ ����#5G��k }��L���� �1CUgy#��$SMON_D�EFPRO ������ *SYSTEM*  ȏ�RECALL ?�}� ( �}�-xcopy f�r:\*.* v�irt:\tmp�back�=>p�ortuc:18700 "	$/-/,?/N+}.�a���0 /�/�/�/Y%0��md:manu�tention.{tpp%emp\,��/$?6?H?[#2�s�:orderfil.datp,,?Ц?�?�?]!)�$b: m/,�?O/OAOT*� t//O�O�O�O_/pO �/�O&_8_J_]?o?�? _�_�_�_�?�?�?�_ "o4oFoYO�O�O�O�o �o�o�O�Ozo_0 B�/�/�/?�����k/buouvrepinceu�i��#�5�G��d*buprog1��n����� ǏZ_l_�_�o!�3�E� �_�_�_�����ßVo ho�o�o�/�A��o�o ��
������ҏ��� ���+�=�P�b����� �����Ϳ��s���� '�9�K�^�ￂ�ϥ� ����ܯ�w���#�5� G�Z�l�~�ߡ߳��� ؿk�}���1�C�Vπh��ߌϝ����T�
�xyzrate 61 m���"�4��F�Y����3192 ���������U���1k�}��� 2D Wiu�������[�9bn�rautou��-?��  �����Z�� |�/1/C/�������/�/�/�/���2317y/�/?.?@? Sev�'?�?�?�? ��v?�(O-O?OR d O�(O�O�O�O�� ��v��#�O&_8_J_]߀�O�;_�_�_�_�6��$SNPX_AS�G 1������Q� P�� '%R[?1]@1.1�_i?��3%oDo'oho Ko]o�o�o�o�o�o�o �o�o.8dG� k}������ ��N�1�X���g��� ����ޏ������8� �-�n�Q�x�����ȟ ��������4��X� ;�M���q���į��� ˯ݯ��(�T�7�x� [�m��������ǿ� ���>�!�H�t�WϘ� {ύ��ϱ������(� ��^�A�hߔ�w߸� �߭�������$��H� +�=�~�a������ ��������D�'�h� K�]������������� ����.8dG� k}����� �N1X�g� �����/�8/ /-/n/Q/x/�/�/�/ �/�/�/�/?4??X? ;?M?�?q?�?�?�?�? �?�?OO(OTO7OxO [OmO�O�O�O�O�D�T�PARAM ���U�Q �	U��JPXTXP�X�OFT_KB_CFG  %S�U?T�PIN_SIM  �[4V�_�_�_�7P�PRVQSTP/_DSBn^4R�_|"X�@SR �qY � & �_�/o%P<VTHI_�CHANGE  �%T\WOaG�RPNUMOV �djOP_ON_E�RRYhZY�aPTN� qUc`�AKbRING_�PRy`�n�@VD�Tsa 1�Ya`  	8W"X0 BTfx���� �����,�>�P� b�t���������Ώ�� ���(�:�a�^�p� ��������ʟܟ� � '�$�6�H�Z�l�~��� ����Ư����� � 2�D�V�h�z������� ¿Կ���
��.�@� R�y�vψϚϬϾ��� ������?�<�N�`� r߄ߖߨߺ������ ��&�8�J�\�n�� �������������� "�4�F�X�j������� ����������0 WTfx���� ���,>P bt�������?SVPRG_CO7UNTOV��a^UN"ENB�o	%M3#�|eA/UPD 1�>kT  
�%R �/�/�/�/�/�/�/? ?,?>?g?b?t?�?�? �?�?�?�?�?OO?O :OLO^O�O�O�O�O�O �O�O�O__$_6___ Z_l_~_�_�_�_�_�_ �_�_o7o2oDoVoo zo�o�o�o�o�o�o 
.WRdv� �������/� *�<�N�w�r������� ��̏ޏ���&�O� J�\�n���������ߟ�ڟ���'�"�4� +Y?SDEBUG y ��J�da)l�SP_�PASS%B?~~�LOG �x%+c#J�G�T��  �]!J�
M�C:\��Z���_M�PC��x%,�>�x!��\� x!�SAV ѳ�Ф�J���SV_�TE�M_TIME 1U�x)��(Ѡ�ͤ��G���T1SV�GUNSs %'�a%�	�ASK_OPTION x%]!:'!)�_DI��4/�E�BCCFG �л�� ���ό�`����������� ���7�"�[�F��j� �ߵߠ���������!� �E�0�B�{�f������������J� 	�8�
�k�}���Z��� ��������c�;��� #I7m[�� �����3! WE{i���� ���//-///A/ w/](H��/�/�/�/�/ ]/?�/?9?'?]?o? �?O?�?�?�?�?�?�? �?�?OGO5OkOYO�O }O�O�O�O�O�O_�O 1__U_C_e_g_y_�_ �_�_�/�_�_o-o?o �_coQoso�o�o�o�o �o�o�o)M; ]_q����� ���#�I�7�m�[� �������ŏǏُ� ��3��_K�]�{����� �ß��ӟ����/� A��e�S���w����� ����ѯ���+��O� =�s�a�������Ϳ�� �߿��%�'�9�o� ]ϓ�I��Ͻ������� }�#��3�Y�G�}ߏ� ��o��߳�������� ��1�g�U��y�� ��������	���-�� Q�?�u�c��������� ������;M_ ���q����� �%I7m[ }�����/ �3/!/C/i/W/�/{/ �/�/�/�/�/�/�//? ?S?	k?}?�?�?�? =?�?�?�?OO=OOO aO/O�OsO�O�O�O�O �O�O�O'__K_9_o_ ]_�_�_�_�_�_�_�_ o�_5o#oEoGoYo�o }o�oi?�o�o�o �oC1Syg��v��p�$TBCSG_GRP 2Շu��  ��q 
 ?�  �����@� *�<�v�`������r�s���|d0�ہ?�q	 HD;)̪�&ff������B\�r�!��333?���!�#�툇L�͇�L�����Cw����ϖ~��CA�C4����Ř@�� ����Ř$���HA���@�p�� ����¯�����
�կ��5�R�a�7�p  �,	V3.0�0�r	r2d7a�	*�����r��hk���(�p7� �\���  ������M�&�-ÿqJCFoG هu�q��-��W���-ς���Ϩ϶� �p������ ���$�� H�3�l�W�iߢߍ��� ����������D�/� h�S��w������ ��
���.��R�d��r �`o�����=������� ���� D/hz ��Y����� �q�A�QSe ������/� /=/+/a/O/�/s/�/ �/�/�/�/?�/'?? K?9?o?]??�?�?�? �?�?�?�oO)O�?IO kOYO�O}O�O�O�O�O �O__1_�OA_C_U_ �_y_�_�_�_�_�_	o �_-oo=o?oQo�ouo �o�o�o�o�o�o) M;q_��� ������7�%� [�I�k���;O����͏ w������!�W�E� {�i�����ß՟���� ���-�S�e�w�1� ������ѯ������ �)�+�=�s�a����� ����߿Ϳ���9� '�]�Kρ�oϑϓϥ� ��������#�5�ߏM� _��ߡߏ��߳��� �������C�U�g�%� w����������	� ���?�-�c�Q�s��� ������������ )_M�q�� ����%I 7m[}��A� ��/�3/!/C/i/ W/�/{/�/�/�/�/�/ ?�//??S?A?c?�? �?�?g?y?�?�?O�? +OOOO=O_O�OsO�O �O�O�O�O�O___ K_9_o_]_�_�_�_�_ �_�_�_o�_5o#oYo ko/�o�o/Qo�o�o �o�o/UCy ��[m���� �-�?�Q��u�c��� ����Ϗ������ ;�)�K�q�_������� ��ݟ˟���7�%� [�I��m�������ٯ ǯ��wo�o'�9��� W�i�����ÿ���տ ��/�A���e�S�u� wωϿ������ϯ�� �=�+�a�O�q�s߅� �ߩ��������'�� 7�]�K��o����� ��������#��G�5� k�Y�����K������� ����1ACU �y�����	��-Q;  w{ {�{��$TBJOP_�GRP 2�C��  K?�{	��ܵ��K� �`pp�� ���� � � {� @w�	 ��D)�+%C2
C랔{�G"�333O!>����K/! LY p$<���d+!? !p$B` w A�A$������'+/=/O%O"�/�*<�+�~-C  B�{@!/?�/�/pF'p%�%p=���5<ҙ*"P!p!��Cz!0�$�?�;C��6���Cуp��.�?K�%p ;��:CAৃ"P$C�C4�?VO�?��?m(�Oj;(A�=�/JhAH�0 YO�OiO�{O_+^fff?U<:f�/F !�0?B�@ f_x_+_�_�Y�_�_�_ �_o�_�_!o;o%o3o ao�omo'o�o�o�o�o��o"�D�{�  ��G%	V3.00��r2d7��*mp�v{�w �GO �~d�� G�0G�� G��| G�: G��� G�� G��t G�2 G��� Gݮ G��l G�* G��� HS�rF�j` �~� F��q � GX �G/� GG8 �G^� Gv �G�ĺs�4 G��� G�� G��\ G� =^p =#�
|8(1DCq�j�k�}�{��?�X�����ESTPAR�p�o��HRրAB_LE 1ݵ��{���� ��v��������z���	���
�����{��������RDI����!�3�E�W�i�єOٟ��� ��+�=��Sן� �����"�4�F�X� j�|�������Ŀֿ� ����0�B�TϚ֠ گ	���~�������`��r����������{�N�UM  C*� � �̐��_CFG ��d��!@�IMEBF_TT܁ս逦�VERʓ���ֽ��R 1ߵ' 8x{v� F��  ��%� 7�I�[�m����� ���������!�3�E� ��i�{����������������_b̐/ �?  k�����T��6����9��I��/ �LTA_�6����L�6���B���/ 7�����/ 
��:���);^��gp]o  ��R�ƙs/ Vudà��/ W�����
�/ [?X�s%�	/����_^���@���ӀMI_CHAN�� �� �#DBGLVL����ҁ� �ETHERAD �?��� ���������/?ˈ� RO�UT��!��!�54S?&<SNMAS�K�(���!255.�5Ys�?�?�?YsӀ�OOLOFS_D�I�pM%�)ORQCTRL �������1NT OUOgO yO�O�O�O�O�O�O�O 	__-_?_Q_c_u_�\�O�_�_�_ЃPE_�DETAI�(�:P�GL_CONFI�G �d�tф��/cell/$�CID$/grp1�_FoXojo|o�oD��?�o�o�o�o �o7I[m�  �������� E�W�i�{�����.�Ï Տ�������A�S� e�w�����*�<�џ� ����+���}��a� s���������)ѽ_�­����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� Ϥ϶��������ύ� "�4�F�X�j�|�ߠ� ������������0� B�T�f�x������ ���������,�>�P� b�t�����'������� ����:L^p ��#���� �$`�EUs�er View �4oXjI�}1234567890� ������@ c/��;2q=/O/ J�s/�/�/�/�/�/=�//C3�/!?3?b/ W?i?{?�?�?�?�/�/<4�?OOF?;OMO�_OqO�O�O�?�?<5 �O�O�O*O_1_C_U_ g_y_�O�O<6�_�_ �__oo'o9oKo]o�_�_<7eo�o�o�_ �o�o/Apo�o<8I���o������%�TF� ��ECameraFx�������� ҏ�����E��9� K����x��������� ҟ�`�+/�'���K� ]�o��������ɯۯ �8��#�5�G�Y�k� 2�pu`�?��ÿ�� ����/�Aϸ�e�w� ��Կ�Ͽ�������� ~����?M�_ߞσߕ� �߹�����T���%� p�I�[�m����� ���O����:��1�C� U�g�y��ߝ������ ����	-?� �_�������� ��9K]�� �����R���o !/3/rW/i/{/�/�/ �/(�/�/�/D/?/? A?S?e?w?�����? �??�?OO)O;OMO �/qO�O�O�?�O�O�O �O__�?��9!_Z_ l_�O�_�_�_�_�_�_ aOo o2o}_Vohozo��o�o�o'_qt	a�0 �o�o	Ho-?Qc u��_�������)�;�M��o�l1 Y������ɏۏ��� �#��G�Y�k����������şן�`��l2 ��/�A���e�w����� ����6�����R�+��=�O�a�s������l3 ��˿ݿ���%�7� I�[�үϑϣ���π�������!ߘ��l4 -�g�y߸ϝ߯����� ����n��-�?��c�u�����4��l5 ����T�9�K�]�o� ����
������&����#5GY���l6 e������� /��Sew��������lz  w	+/=/O/a/ s/�/�/�/�/�/�/�+   /	/'?9? K?]?o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_	o�o-o?oQoco�,  }
s (  � ( 	 so�o�o �o�o�o�o%'�9o]���}j: �K�� � �D�V�h�z�����u �ȏڏ�3��"�4� F�X�j����������� ֟�����0�w�T� f�x���������ү� ��=�O�,�>�P���t� ��������ο��� �]�:�L�^�pςϔ� ۿ������#� ��$� 6�H�Zߡϳϐߢߴ� ��������� �2�y� V�h�z��ߞ������ ����?��.�@���d� v������������� _�<N`r� ������% &8J\���� �����/"/i {X/j/|/��/�/�/ �/�/�/A/?0?B?�/ f?x?�?�?�?�??�? �?OO?,O>OPObOtO8�O�?�p@ �B�O��O�O�C�G�`����O_&_8_J_\_n_ �_�_�_�_�_�_�]_ o o2oDoVohozo�o �o�o�o�o�o�_
 .@Rdv��� ����o��*�<� N�`�r���������̏ ޏ���&�8�J�\� n���������ȟڟ� ���"�4�F�X�j�|� ������į֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tφϘϪϼ�t���I(A �O��$TPGL_O�UTPUT �|�1�1 ���,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p�������������  �2345678901����%�7�I� Q��2��x��������� ��j���,>P��}Z����� bt $6HZ �h�����p �/ /2/D/V/� / �/�/�/�/�/�/~/�/ ?.?@?R?d?�/r?�? �?�?�?�?z?�?O*O <ONO`OrO
O�O�O�O �O�O�O�O�O&_8_J_ \_n___�_�_�_�_ �_�_�_o4oFoXojo |oo�o�o�o�o�o�o�o��}��0BTfx��}@�Ͽ���>��( 	 ��� �*��N�<�r�`��� ����̏����ޏ�� 8�&�H�n�\������� ��ڟȟ����4�"��X���OFF_L�IM#��������t�N_SV�x�  ����P_MON ������������STRTCHK ���-��VTCO�MPAT��)���VWVAR 뿭�"�N���  � �d���Ң�_D�EFPROG �%�%
OUVR�EPINCE  ���AUTO{���ISPLAY#���INST_MSK�  � кI�NUSER�ִL�CK(��QUIC�KMENL�ִSC�REk��*�tpscִ(���h�Ɋ���_��ST����RACE_CF�G ��L��Ϡ	��
?����H_NL 2�L��S� y�?�Q�c�u���ߙ߽߫�����IT�EM 2�+� �%$�  =�<�B�T�\�  !b�j�v�&� ���4����j���� ��i���������@� 0�B�T�n�x�����H n����,� P�"4�@�� �d���L� p�K/�f/��/�/  /�/$/v/�/Z/?~/ *?P?b?�/n?�/�/? �?2?�?OOz?:O�? �?�?FO^O�?�O�O.O �OROdO-_�OH_�Ol_ ~_�O�___�_<_�_ `_o2o�_�_�_�_�_ �_joo�o�o�o\o �o�o�o�ot�� �4FX�*�� N�`��l���Ï� ޏB���x�*���� w�ҏ������ȟڟ>� �b�t��� ���V�|� ��򟲯�(�:���֯ p�0�B���N�ʯܯ��  ���$����Z��~�(��Y���S�����^ʟ�  ��^�q ѵ���
 ��������d�R_GR�P 1���� 	 @��L�^ۀH�~�lߢߐ��ߴޠ ���������%��I�4�?�  d�v�`� ������������� �8�&�\�J���n���������	,��� ~)�SCB 2�z� O�L^p�������d�X_�SCREEN 1��7�
 �}i�pnl/gen.htm�<N`�r�&�Pan�el setup�}������/"/ ��Z/l/~/ �/�/�/+/�/O/�/?  ?2?D?V?�/�/�?�? �?�?�?�?]?�?�?.O @OROdOvO�O�?�O#O �O�O�O__*_�O�O `_r_�_�_�_�_1___ U_oo&o8oJo\o�_ �o�_�o�o�o�o�o�o�uo�UALRM_�MSG ?7���� _zQc� ���������6�)�Z�M�~�2uSEoV  @}��0rEt��zϭ���}A��   B������7��%�7�I� [�m��������ǟ՗4��1��Ƌ ?�4�����A��*SY�STEM*&�V8�.1079 G�1�/30/2013� A 7��5�"��UI_MENH�IS_T   �8 $q�T_H�EAD��}�EN�TRY ��$�DUMMY2 k ��3��  j��OUSEt���$ACTION���$BUTTˤR�OW͢COLUM�̣TIME��$�RESERVED���j�PANED�ATt� � �$PAGEURL� }$FRA��)$HEL�P�PA'�TER�1+�<���H���H�4�F�5F�6F�7F�86+�INB�VA ����	�STAT*���1xr����� j�USRVIEWt�� <Ġn�U!���NFIG��FO�CUS��PRIM�!�m�����TRI�PL*�m�UND�O_t�t�  �$4�ENB��$WARNJų���__INFOt�y���_PROG �%$TASK_�I��t�OSIDX҈�R��`�TO�OLt� 4 �$X��$����Z\��ߡ$P��R��F��NU�9`�U&�Bt��������E���`�OFF��u� �D{���O?� 1���)�Q���GU�N_WIDTH � ��K�_SU�B��  
`�R�T���t�	��$qD����ORN�ׯRAUX��T��E�NAB-���VCC�M��� 
$�VISʠ_TYP�ɳC(�RA��PO�RTХ�A�C���N^(�%$EX��_��$��_F�P��P�� A��a�LU ��$OUTPUT_�BM�
���MR�_���h �����+�DRIV�����SET_VT�C���BUG_C�ODɴMY_UB	Yȴ6�	����ʠE���,���:�f�x�O�HANDEY��E�8p�ULX�P��AL_����GD_SPA�CIN���RGT ������������U�RE����U��w��������  6��RG��PNT�r��R���� dġ�Xr�FLA���	�T�AXS���SW���_A��y���S���O�BA��zy�	$E��UE���yз���HK��r �
�MAXv{ER��MEAN�	�WOR��z��MR�CV�� ��O�RG9pT_C&�P )�
REF ���-�i ����N�b b18��_RC��@�� 8���M���M����� ��P�űG]����$GROUP����:&��� ��;2p CREǰw�.�$�Ab"N!�HK��SULT����COVE��Y��a NT6��%����&���&ձ�#m L�6��%F��%���'ձ����9�0 m&z#PAu� z#oCACHO�LOV�*4@1��E9���C�_LIMIf3FR�n8TDn8�$HOt��=�.0COM������OBO�8(� |�!$IN_VP��<���2_SZ3�#�56�#�512���8R���:TKQ�8o0�8W�A5MPBJFAIjo0G�?0ADrI�U�IMRE $�B_�SIZ/$PM��N�D� P�ASYNB{UFP�VRTD�E��D�A�3OLE_2�D_��EW�PC&��TUq�@0Q� �E�ECCU��VEM���)54Ro6 ��$���� CKLAS�v�	�VLEXEJ5G��� �z!nO�FLDd�DE�C�FI�@�W� �W���V;�s� (����UF�QǠ��! ��_��L�#���Q�� hP �1���!��K�$��$�=�E�!}�C�U�%$"A7
�@PS�Kt4M:&�e  ���TRbUt�� $p TIT-���A0=�OPɤ��VSHIF:��`��|!#����URO�d _R�@�+t H�C=u��L�^�p�o0`���qi �ҏsTI�!N�tSCO'r�sC�� ��S¨�SwS£vS� �wS¾x����Ꞣ���s�ED���w� m SM7�A��$ADJ�`K�%�UA_{"u�A��g�}�LIN.����ZABC������
��ZMPCF���  C��J���LN�`�a��I��� ���1� ���CMCM��C�3COART_6��Pa? $JT�N�D�1Z�k�d���p���ΎUXW����UX!E�񞖙�_���u����������ɖ߁PB5��r�������uY��Dc� y�:2v/�IGH���h#?(p ���$  � �d7ۀK$Bm KK�]a_�b,�#u�RVn0F��cOVC��O�D��$P�`��Ǳǡ
�Iݣ��5D�TRACE�J�Va��SPHE}R�� ! ,p �1�G�Y��$�DE�Fx�?%����c��^�(%�ހx���t����� ѿ�������*�O��:�s�^ϗϢ�T�IN.��  c��Ϧϵ_T`H��1 c���(��� ��(/SOF�T͡/GEN��K�?current�=menupage,153,1��pT�f�xߊ߀� �.�962A�������0�߭߿�36��Z� l�~��������� ������7�I�[�m� ��� ����������� ��3EWi{� �.����'��ѶSew �������/ /+/�O/a/s/�/�/ �/8/J/�/�/??'? 9?�/]?o?�?�?�?�? F?�?�?�?O#O5O�? �?kO}O�O�O�O�OTO �O�O__1_C_.@ y_�_�_�_�_�_�O�_ 	oo-o?oQo�_uo�o �o�o�o�o�opo );M_�o��� ���l��%�7� I�[�m��������Ǐ ُ�z��!�3�E�W� i�T_f_����ß՟� �����/�A�S�e�w� �������ѯ���� ��+�=�O�a�s���� ����Ϳ߿�ϒ�'� 9�K�]�oρϓ�"Ϸ� ��������ߠ�5�G� Y�k�}ߏ�z������� ������"�C�U�g� y���,�>������� 	��-���Q�c�u��� ����:������� )����_q��� �H��%7 �[m��������$UI_PA�NEDATA 1������  	�}��/ /2/D/V/h/ )j/�/�$��/�/�/ �/??z/7??[?m? T?�?x?�?�?�?�?�?�O�?3OEO,OiOvI� ���B�/�O�O �O�O�O _SO$_�/6_ Z_l_~_�_�_�__�_ �_�_�_o2ooVo=o zo�oso�o�o�o�o�o
}L+v�H_M_ q����o�>_� ��%�7�I��m�� f�����Ǐُ����� !��E�W�>�{�b��� ��$6�����/� A���e���������� ѯ���\�� �=�$� a�s�Z���~���Ϳ�� �ؿ�'��KϾ�П �ϓϥϷ�����.��� ߄�5�G�Y�k�}ߏ� �ϳߚ���������� 1�C�*�g�N���� �����X�j�(�-�?� Q�c�u��������� ����)��M_ F�j����� �%7[B �������/ !/tE/��i/{/�/�/ �/�/�/</�/�/?? A?S?:?w?^?�?�?�? �?�?�?O�?+O�� aOsO�O�O�O�OO�O �Od/_'_9_K_]_o_ �O�_z_�_�_�_�_�_ o#o
oGo.oko}odo`�o�o�o8OJO}��o@!3EWi)�o �U}����� �{8��\�C�U��� y�����ڏ�ӏ����4�F�-�j�v�TCNK��$UI_POST�YPE  TE�� 	 �v�͟��QUICK�MEN  �����П��RESTO�RE 1TE�  � ]�G�A�S�w�mr��� ����ѯ㯆���+� =�O��s��������� f�ȿڿ�^�'�9�K� ]�o�ϓϥϷ����� �ϐ��#�5�G�Y�� f�xߊ����������� ��1�C�U�g�y�� ���������ߚ�� ���:�c�u������� N���������; M_q�.���� &�%7�[ m���X����/!/ۗSCRE��?�uw1sc<�u2\$U3\$4\$5\$6\$�7\$8\!��USE�R> C/U"T= ^#k�sf#�$4�$5�$6��$7�$8�!��ND�O_CFG ��`�a��PDAT�E �)��Noneޒ� _I_NFO 1�&Q0��0%'/l?x8Z?�? ~?�?�?�?�?O�?+O OOOaODO�O�OzO�O�Ԝ>1OFFSET ��OS5� �__0_B_o_f_x_ �_�_�_�O�_�_�_o 5o,o>okoboto�o�[� ��m
�o�o�HUFRAME  �d�6;1RTOL_�ABRT932rE�NB;,xGRP �1	0���Cz  A��s�q�a������v��*z��U[x1J{MSKG  ^uQ3LyNq�%I:%�o��ݒV�CCM_PAp �
<%~�VSCAM1 *Xߏ焣����5�����MRwr2���Ҁ�?��	с��	`ֆ�Z�1B��5��A@�pp�pȣ� �o��������@�<������u�A���T�Z�? B���o�Z� s�����۟����ܯǯ  ��$��!�Z���;� ��{���ƿy�������ISIONTMOiU:p^�˅����"f`��f�`�@�q F�R:\�\0A\�� �� M�CT�LOGa�  � UD1T�EX��ϰ�' B@ �������������� ��  =	 1-� n6  -�� t������, ֌�_�=�̩�h����z�TRAIN��$�4��� (��h��� �����������"�4� j�X�n�|������^��LEXE<���11-80��MPH?ASE  &53yk���R 2�
 ��]�o��������a������ ���� $6*1�l��������� ����s����������G	n�opqr�stuvw Z�~�� �����./f </n`/r/��/�/�/�/�//h$/?H/ &?L?~/p?�?�?�?�? �?/? O2?$O6Oh?�ZOlO~O�O�OD��u�3� �?�OO__LO>_P_�b_t_�_D��D	��BH
�O�_�O �_o4_&o8oJo\ono�H�@~		�3�?
�
��Æ�o �_�o�oo&8�J|o�3�
�
g�hijk �@\��o��o�o����&�8�ƃ��SH�IFTMENU Y1>�c�<��%����&���t���ӏ�� ��	����?��(�N� ��^�p��������ʟ ܟ�;��$�q�H�Z�0��~�T��[�K���	VSFT1���~VSCAM�5ذ?��!�@z`��G�  A�ٰU8ٰٰ��p*��$���"�!����s�L�̦MEP �la�/� T�MO����zR�WAITDINEND �� �w���OK  �Oյ��ԿS迻�T�IM����G ��5�ǿX��8��8�<%Ϲ�RELE9�h��s���TM��s��~��_ACTIV���1ѹ�_DATA [�2�%��h�,���RDISg�����$ZABC_G_RP 1۩I��,�qp�2p�t�ZMPCF_G 1�v��I�0�������M�P��۩/��'�q���'�s�8��`���_����?��� �����/����V�������`�[��������������Ѕ������P_CYLINDER 2��� Н� ,(  *m~��j���� �� %gH�lSe� ����-/�� D/+/h/O/��/�/���=�2 ۧ4� � ��/<�~�3??W?�e:�/�?�7��1A��;SPHERE 2!M�/�?R/�? O�?8O�/�?nO�O� �OCO)O�O�O�O�OWO 4_F_�O�O|_�O�_�_��_�__�_oo��ZZ�� ���