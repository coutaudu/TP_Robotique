��   D�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A 
  ����CELLSET�_T   �w$GI_STY�SEL_P }7T  7ISO:iRibDiTRA�R�>�I_INI; �����bU9AR�TaRSRPNS�1Q234�5678�Q
TROBQACKSNO� �)�7�E�S �a�o�zU2 3 4 5 6 7 8awn&GINm'D�&��) %��)4%��)P%�̖)l%SN�{(OU���!7� OPTNAA�73�73.:B<;�}a6.:C<;CK;C�aI_DECSN�A�3R�3�TRY�1��4��4�PTHCN�8D�D�INCYC@HG��KD�TASKOK �{D�{D�7:�E� U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V�8�Tb@SEGq�Tp��T�@REQ� d�drG�:Mf�GJO_HFAUL�Xpd�dvgALE�  �g�c�g�cvgE� �H<�dvgNDBR�H�dgRGAB�Xtb�	  �CLML�Iy@   �$TYPESI�NDEXS�$$�CLASS  O���lq�����apVIRTUA�Li{q'61ION�  ��c��q�t+ UP0 ��u�qSty�le Select 	  ��r�u�Req. /Ec�ho���yAck����sInitGiat�p�r�s�t@�O�a�p���;pV �����������q����𱇪q��sOpti�on bit AJ��B����C��Decis�co�d;��zTryou�t mL��Pat�h segJ�nt�in.�II�yc�:��Task O�K��!�Manual opt.r�pIAԖBޟԖC�� decsn ِ��Robot i?nterlo�"�>>� isol3���C��i/�"�z�ment��z�ِ����~_�status��	MH Faul�t:��ߧAler���%��p@r 1�z L��[�m�+��; LE_COMN�T ?�y�   ��䆳�Ŀֿ� ����0�B�T�g�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼�������������U������   ���ENAB  ���u�����x���ꐵMENU>���y��NAME ?=%��(%$*4��� D��p2�k�V���z��� ����������1 U@Rdv��� ����*< u`������ ��/;/&/_/J/f/ n/�/�/�/�/�/?�/ %??"?4?F?X?j?�? �?�?�?�?�?�?�=