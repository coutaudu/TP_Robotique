��  Ij�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����SBR_T �  | 	$SV�MTR_ID � $ROBOT�9$GRP_�NUM<AXIS�Q6K 6NFF~3 _PARAMF�	$�  �,$MD SPD_[LIT  &2*�� � �����$$CLASS ? ���������� VIRT�UAL��'  1� � T����R-20�00iB/165�F��:AC�aiSR 3' �80A��
H1� DSP1-S1���	P02.0�29,  	�  ��P�aR� �# ��w������ ���
=�#�2r�9  ~���%����8� l� � ����?� ��� ץ���< �""��������	  �3�4��<�����ow����������� ( 	���� �����O��������	 ������_�����qc�9	`B 0� ��� ��� :?�p�:@  ?'bx�E/�/0�/�/�/���/?�3?C?U?��Z����5'h���;��|����j�6��\��:'�����L"-#\?�?�h0	BT2^qj|���	��U����^p��@��� ���������- 4�k�
 x�Y��W}���qs+��, %� ��4 �8$Q|�?����S\'o��;j/ �~/ �/�!:@�/r_�_�_�_�?�_'?�_o]?o? �6��0����/��V�6%�0�����k�"��oso��$�?0�?T3^�RP"O4K��GKp���^tO�x�BC�G9 �3F30���^% +����=����0���D���� ��/�� W8$ozo�������\'��a"_ �6_H_Z_ #�5�G�Y��_}��_�� ��ŏ o�����1�qab�o4�b/12/4N4SY�4^4�o�lc:~�e�q����2�P��{Pu���t�k0���n$(H���@���z��Sx.�.�!BA5@#�5���I ���� r8$��E��������\!�E�����EB����  ����o���"��y/m���� 	��v�?��fF�k��}�������ſ׿�I�F�0j�|�5^�5�������>Ɨ���ҟ���
e��;�:�:���������?0 �\�m�8$���z���^��;����p�������ʯ�ߥ߷� ��$���H���#�5�G�`Y�k�}������R0"�|�6^6F��X�j���Ɩ���؊Ϝ���^��=U�0�0��ϛ������KX���� �n8$7$F/��4����}����^�p߂�K]o� �ߥ �����#5GY�����Z�nnJ��	��� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?2<�2?V? h?z?�?�?�?�?�?�? �?
OC�~(O�� ��O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_@?oo ,o>oPoboto�o�o�o �oOJO<O`OrO: L^p����� �� ��$�6�H�Z� l�~����_��Ə؏� ��� �2�D�V�h�z� �o����0��
� �.�@�R�d�v����� ����Я�����*� <�N���r��������� ̿޿���&�8ϴ� ��P�ʟܟ����� �����"�4�F�X�j� |ߎߠ߲��������� �h�0�B�T�f�x�� ���������@�r�d� -��Ϛ�b�t������� ��������(: L^p����� �� $6HZ l~������4� F�X� /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?��? �?�?�?�?�?OO*O <ONO`O��xO�/ /�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4o�?Xojo |o�o�o�o�o�o�o�o hO�O�OU�O�O� �������� ,�>�P�b�t������� ��Ώ��<o��(�:� L�^�p���������ʟ &��\n�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψ�� �����,�>���*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \︿��������� �����"�4����ϴ� }����ϲ��������� 0BTfx� ������d� >Pbt��� ����N�/
/�� ����p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?"�? �?O O2ODOVOhOzO �O�O�O,//�OB/T/ f/._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�?�o�o �o�o�o&8J \�O�O�O� __� ���"�4�F�X�j� |�������ď֏��� ��0��oB�f�x��� ������ҟ����� v?�2�������� ��ί����(�:� L�^�p���������ʿ ܿ�J��$�6�H�Z� l�~ϐϢϴ�����T� F���j�|���V�h�z� �ߞ߰���������
� �.�@�R�d�v��� �����������*� <�N�`�r������� ��(�:�&8J \n������ ��"4FX�� j������� //0/B/��g/Z/�� �����/�/�/�/?? ,?>?P?b?t?�?�?�? �?�?�?�?OOr:O LO^OpO�O�O�O�O�O �O�O _|/n/_�/�/ �/~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�o�o�o0O�o
 .@Rdv�� �_:_,_�P_b_*� <�N�`�r��������� ̏ޏ����&�8�J� \�n����o����ȟڟ ����"�4�F�X�j� ������� ���� ��0�B�T�f�x��� ������ҿ����� ,�>Ϛ�b�tφϘϪ� ����������(ߤ� ��@ߺ�̯ޯ�߸��� ���� ��$�6�H�Z� l�~���������� ��X� �2�D�V�h�z� ����������0�b�T� xߊ�Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/���/�/$ 6H?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfO��O �O�O�O�O�O�O__ ,_>_P_�/�/h_�/�/ ?�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $�OHZ l~������ �X_�_|_E��_�_z� ������ԏ���
� �.�@�R�d�v����� ����П,���*� <�N�`�r��������� �߯үL�^�p�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώ�ꟲ��������� ��0�B�T�f�x��� 毐�
��.����� ,�>�P�b�t���� ����������(�:� L���p����������� ���� $�߲ߤ� m���ߢ���� � 2DVhz �������T� 
/./@/R/d/v/�/�/ �/�/�/�/>?�/t ��`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O/�O �O�O_"_4_F_X_j_ |_�_�_??�_2?D? V?o0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt�O�� ������(�:� L��_�_�_���_oʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �|2�V�h�z� ������¯ԯ���
� f�/�"����������� ����п�����*� <�N�`�rτϖϨϺ� ����:���&�8�J� \�n߀ߒߤ߶���D� 6���Z�l�~�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt����� ��*��(: L^p����� �� //$/6/H/�� Z/~/�/�/�/�/�/�/ �/? ?2?�W?J?� ���?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O_b/*_ <_N_`_r_�_�_�_�_ �_�_�_l?^?o�?�? �?no�o�o�o�o�o�o �o�o"4FXj |���� _�� ��0�B�T�f�x��� ���_*oo�@oRo� ,�>�P�b�t������� ��Ο�����(�:� L�^�p��������ʯ ܯ� ��$�6�H�Z� ���r�����ؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.ߊ�R�d�v߈ߚ� �߾�������� ��0謹��ο���� ��������&�8�J� \�n������������� ��H�"4FXj |���� �R�D� h�z�BTfx� ������// ,/>/P/b/t/�/�/�� �/�/�/�/??(?:? L?^?p?�?��?�? &8 OO$O6OHOZO lO~O�O�O�O�O�O�O �O_ _2_D_V_�/z_ �_�_�_�_�_�_�_
o o.o@o�?�?Xo�?�? �?�o�o�o�o* <N`r���� �����p_8�J� \�n���������ȏڏ �Hozolo5��o�oj� |�������ğ֟��� ��0�B�T�f�x��� �������ү���� ,�>�P�b�t������� �Ͽ¿<�N�`�(�:� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~�گ�ߴ������� ��� �2�D�V�h�� ֿ����������
� �.�@�R�d�v����� ����������* <��`r���� ���p��� ]�������� ��/"/4/F/X/j/ |/�/�/�/�/�/�/D �/?0?B?T?f?x?�? �?�?�?�?.�?�?d v�PObOtO�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_?�_ �_�_ oo$o6oHoZo lo~o�oO�?�o"O4O FO 2DVhz �������
� �.�@�R�d��_���� ����Џ����*� <��o�o�o���o�o�� ̟ޟ���&�8�J� \�n���������ȯگ ����l�"�F�X�j� |�������Ŀֿ��� V��ό�����xϊ� �Ϯ����������� ,�>�P�b�t߆ߘߪ� ����*�����(�:� L�^�p�����4� &���J�\�n�6�H�Z� l�~������������� �� 2DVhz ��߰����
 .@Rd������ �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?� J?n?�?�?�?�?�?�? �?�?O"O~GO:O� ���O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_R?o ,o>oPoboto�o�o�o �o�o�o\ONO�orO�O �O^p����� �� ��$�6�H�Z� l�~�������o؏� ��� �2�D�V�h�z� ���o՟0B
� �.�@�R�d�v����� ����Я�����*� <�N�`���r������� ̿޿���&�8�J� ��o�b�ܟ� ����� �����"�4�F�X�j� |ߎߠ߲��������� ��z�B�T�f�x�� �������������� v� ��ϬϾφ����� ��������(: L^p����� �8� $6HZ l~����B�4� �X�j�2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?� �?�?�?�?�?OO*O <ONO`OrO��O�O/ /(/�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFo�?jo |o�o�o�o�o�o�o�o 0�O�OH�O�O �O������� ,�>�P�b�t������� ��Ώ����`o(�:� L�^�p���������ʟ ܟ8j\%���Z� l�~�������Ưد� ��� �2�D�V�h�z� �������¿���
� �.�@�R�d�vψϚ� ���ϲ�,�>�P��*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \�n�ʿ�������� �����"�4�F�X��� ��p������������ 0BTfx� ������ ,��Pbt��� ����/`����� M/�����/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?4 �?O O2ODOVOhOzO �O�O�O�O/�O�OT/ f/x/@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�?�o �o�o�o&8J \n��O�O�_$_ 6_��"�4�F�X�j� |�������ď֏��� ��0�B�T��ox��� ������ҟ����� ,����u����� ��ί����(�:� L�^�p���������ʿ ܿ� �\��6�H�Z� l�~ϐϢϴ������� F���|�����h�z� �ߞ߰���������
� �.�@�R�d�v��� ����������*� <�N�`�r�������$� ���:�L�^�&8J \n������ ��"4FXj |������� //0/B/T/������ �/��
�/�/�/?? ,?>?P?b?t?�?�?�? �?�?�?�?OO(O� :O^OpO�O�O�O�O�O �O�O __n/7_*_�/ �/�/�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�o�o�o�oBO
 .@Rdv�� ���L_>_�b_t_ �_N�`�r��������� ̏ޏ����&�8�J� \�n������� ȟڟ ����"�4�F�X�j� |��
��ů �2��� ��0�B�T�f�x��� ������ҿ����� ,�>�PϬ�bφϘϪ� ����������(�:� ��_�R�̯ޯ���� ���� ��$�6�H�Z� l�~���������� ���j�2�D�V�h�z� ��������������t� f��ߜ߮�v�� �����* <N`r���� �(��//&/8/J/ \/n/�/�/�/ 2$ �/HZ"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO� �O�O�O�O�O�O__�,_>_P_b_�%�$S�BR2 1�%��P T0 � �/�) �_�_�_ �_oo&o8oJo\ono �o�o�o�o�_�_�o�o "4FXj|� �����o�o�o� 0�B�T�f�x������� ��ҏ�����,�� P�b�t���������Ο �����(�:��^� A���������ʯܯ�  ��$�6�H�Z�l�O� ��s���ƿؿ����  �2�D�V�h�zόϞ� ��j_��������&� 8�J�\�n߀ߒߤ߶� ���ٸ���
��.�@� R�d�v������� ��������*�<�N�`� r��������������� &
�6\n� ������� "4FX<|�� �����//0/ B/T/f/x/�/n�/�/ �/�/�/??,?>?P? b?t?�?�?�?�?�/�? �?OO(O:OLO^OpO �O�O�O�O�O�O�O�? _$_6_H_Z_l_~_�_ �_�_�_�_�_�_o o _DoVohozo�o�o�o �o�o�o�o
.@ R6ov����� ����*�<�N�`� r���h����̏ޏ�� ��&�8�J�\�n��� ��������ڟ���� "�4�F�X�j�|����� ��į֯�����0� B�T�f�x��������� ҿ�����,�>�P� b�tφϘϪϼ����� ����(�:��^�p� �ߔߦ߸������� � �$�6�H�Z�l�Pߐ� ������������ � 2�D�V�h�z������� ��������
.@ Rdv����� ���*<N` r������� /�&/8/J/\/n/�/ �/�/�/�/�/�/�/? "?4?/X?j?|?�?�? �?�?�?�?�?OO0O BOTO8?J?�O�O�O�O �O�O�O__,_>_P_ b_t_�_jO�_�_�_�_ �_oo(o:oLo^opo �o�o�o�o�_�o�o  $6HZl~� ������o� � 2�D�V�h�z������� ԏ���
�� �@� R�d�v���������П �����*�<�N�2� r���������̯ޯ� ��&�8�J�\�n��� d�����ȿڿ���� "�4�F�X�j�|ώϠ� �ϖ���������0� B�T�f�xߊߜ߮��� ��������,�>�P� b�t��������� �������:�L�^�p� ��������������  $6�Fl~� ������  2DVhL��� ����
//./@/ R/d/v/�/�/~�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�/�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O�? "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o _Tofoxo�o�o�o�o �o�o�o,>P bFo������ ���(�:�L�^�p� ����x��ʏ܏� � �$�6�H�Z�l�~��� ������������ � 2�D�V�h�z������� ¯ԯ�ʟ���.�@� R�d�v���������п �������<�N�`� rτϖϨϺ������� ��&�8�J�.�n߀� �ߤ߶���������� "�4�F�X�j�|�`ߠ� ������������0� B�T�f�x��������� ������,>P bt������ ��(:L^p ������� / /�6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?(/h?z?�?�?�? �?�?�?�?
OO.O@O ROdOH?Z?�O�O�O�O �O�O__*_<_N_`_ r_�_�_zO�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�_�o�o "4FXj|�� ������o�0� B�T�f�x��������� ҏ�����,��P� b�t���������Ο�� ���(�:�L�^�B� ��������ʯܯ� � �$�6�H�Z�l�~��� t���ƿؿ���� � 2�D�V�h�zόϞϰ� �Ϧ�����
��.�@� R�d�v߈ߚ߬߾��� �������*�<�N�`� r����������� ����
�J�\�n��� �������������� "4F*�V|�� �����0 BTfx\��� ���//,/>/P/ b/t/�/�/�/��/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�/ O O$O6OHOZOlO~O�O �O�O�O�O�O�O_�? 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o $_dovo�o�o�o�o�o �o�o*<N` rVo������ ��&�8�J�\�n��� �����ȏڏ���� "�4�F�X�j�|����� ��ğ��������0� B�T�f�x��������� ү���ڟ�,�>�P� b�t���������ο� ���(��L�^�p� �ϔϦϸ������� � �$�6�H�Z�>�~ߐ� �ߴ���������� � 2�D�V�h�z��p߰� ��������
��.�@� R�d�v����������� ����*<N` r������� ��&8J\n� �������/ "/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?8/x?�?�?�?�? �?�?�?OO,O>OPO bOtOX?j?�O�O�O�O �O__(_:_L_^_p_ �_�_�_�O�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�_�o  2DVhz��� ����
��o.�@� R�d�v���������Џ ����*�<�N�