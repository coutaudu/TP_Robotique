��   ��A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ��	��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !� FTP�_CTRL. =@� LOG_8	��CMO>$DN�LD_FILTE�R�SUBDIR�CAP���HOv��NT. 4� �H�9ADDRT�YP� A H� NG#THOG��z +�LS/ D $ROBOTIG �BPEER�� MwASK@MRU~;OMGDEVK%�RCM+ �� $�� ��QwSIZNTIM�$STATUS�_�?MAILS�ERV�LANT�� =$LIN�=�$CLU��f=${TOcQ$CC5&{FR5&ALAR��B�TP�\#VA�Rd(�RDM*�� $DIS��� TCPIo/ >3 $ARP�)o_IPFOW_���F_INF=A~LASS��HO_� INFO�z"TELs P�~���� WO�RD  $A7CCE� LV���OU wORT }�ICEUS 0   �$�#  ���r1���
��
g0VIRTUALo?�1'0 ��5
���F������4�5� �� �=��!y1O����$ETH_F�LTR  �6�3� ���������K�� �=2K�"S�HAR� 1�9�  P O�O�4 �O�O�O_�O*_�ON_ _Z_5_�_�_k_�_�_ �_�_o�_8o�_ono 1o�oUo�oyo�o�o�o �o4�oX|? u������� �*��S�x�;���_� ����䏧��ˏݏ>� �b�%���I���m�� �����ǟ(��L�� E���q���i�ʯGz �_LIST 1�1Mx!1.�0�ӯ���1���2�55.M������5�2
����0�B�T�f�x�3���������̿޿x�4���q�  �2�D�V�x�5r��@���Ϫϼ���x�6�π�a��"�4�F� ����1�K��}0�� Q����= ��1�C��g�y��^�������Q������ ��9�K�]�o�.����������J$� �>�$ �%� �=��5�5	1���9�@@H!�� X��rj3O_tpd���1 �0>y1!KC�0��m	���6�!C�P0����!GCONn03nzOsmon�