��  �\�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A9  �����ABSPOS_�GRP_T  �  $PAR�AM  ����ALRM_R�ECOV1  � $ALMOEkNB��]ONi�I M_IF1 �D $ENAB�LE k LAS{T_^  d�uU�K}MAX� �$LDEBUG�@  
FPCO�UPLED1 �$[PP_PRO?CES0 � �y1��UREQ1� � $SO{FT; T_ID��TOTAL_EQf� $,NO/�PS_SPI_I�NDE��$DX��SCREEN_�NAME ^�SIGNj�|�&PK_FI� �	$THKYޠPANE7 � 	$DUMMY�12� �3�4����ARG_�STR1 � �$TIT�$I��1&�$��$�$5&6&7*&8&9'0''@�%!'�%5'1?'U1I'1S'1]'2h"�GSBN_CFG�1  8 $�CNV_JNT_�* �DATA_C�MNT�!$FL�AGSL*CHE�CK��AT_C�ELLSETUP�  P� HO�ME_IO� }%:3MACROF2�REPRO8�DR�UNCD�i2SM�p5H UTOBAC�KU0 ��	DEVIC#T�Ih�$DFD��ST�0B 3$�INTERVAL��DISP_UNsIT��0_DO�6�ERR�9FR_F�a�INGRE5S�!Y0Q_�3t4�C_WA�4�12JO�FF_� N�3DEL_HLOG�2�jA��2?�1k@�?Q�� ���H X_�D�#	 d �$CARD_EX�IST�$FS?SB_TYPi� �CHKBD_SE��5AGN G� �$SLOT_N�UMZ�APREV�D�G �1_ED�IT1
 � *h1G=H0S?@f�%$EPY$�OPc iAEToE_OK�BUS�oP_CR�A$�4xJVAZ0LACIw�Y1�R�@k �1CO�MMEc@$D�V�QOk@:Y���$QL*OU/R , $�1V1AIB0~ OL#eR"2�CF�D X �$GR� � S!1�$MB_@NFLI�C�3\`
UIRE�s3��AOMqWI�TCHWcAX_NR.0S�=`_;G0� � 
$WARNM'@f��@� sLI? �aNST� �CORN��1FL{TR�eTRAT@0�T�` �0ACC��1�` |�rOR�I�P�CxkRTq0_sSF� �!CHG]I1 [ TT`4u3I*pTY�2Qq�K*2  x ��`� 1�B*HDR��J* ��q2�v3��v4�v5�v6�v7j�v8�v9��QpO�$ <� Mo_o�qh�s1<`O_MO�R. t �0Ev�NG� �0BA� �Qt�Q}��r��@��v�©�P�0����h�`^P/P�2� �p�Jp_R�bLq�@b�J	r	�$�JV�@�CD��m|gv�uMt�P_}0OF� � ; @� RO_����aIT8C��NOM	_�0�1��q3�@���$ ����|hP���mEX�`G�0�� �0"��`�b
$T�FR�J �D3��T�O�3&@U=0�� ���H�2�T1m�E��� �e��f���f��0CPDB�GDE��@�$`PU�3�fc)���AX 1܁dbETAI�3BU�F�F�����! �� ˧�`PI�U��PL�MK�MX����[�FL�SIMQ�S��KEE��PAT�`�!� ������MCU� �$�}1JB�`-�}1DE�C㺋��FɱT�� �7PCHNS_wEMPvr$GA��'��@_y�q3�`1_�FP͔x�TCR�SPEubw�q0�cg�S�!�� V�A���!�����JR!0��SEGF�RApv r�R�T�_LIN�C��PVEF�M������Y ��P��)B��وD )\�}f�e 	�"��	��.0�Z�p�Ql��SIZCuх�d�To�A��ڭ�>	�RSINF��p ����?���ܭ���s�¸�LItx�1��CRC�eFCCC�`�� >�R��mRMAl� R��P� �$�D�d�c2��C��j@TA����0�@��l���EV���jUF��_��Fw�N��� ��f��!�� 2�\������1C���! ����hRG�Ps�
qF��7bg�qD���2g�LEW(���s� �e�>�P��PqR�D� ��&�pou2|��A6N�HANCI�$LG �`-��1�Pd��@�d�a!A?@l���~0R��z�jME��uAk��e3RAs3jAZC�t��T�OEqFCT�q��`F�`m�g�̰�ADI;� q� � l��`��`�`|�H�aS=P�r��AMP��Ҥ�Y8C?�MAE�S����r�I�$_  *�I���CSX�a�!&�p	$JTpT�X��C_ N�@h�IMG?_HEIGH�A�gWID��h�VTE�:�U�0F_A��- �@EXP(�c-%��CU���QU�1� $`TIT�1�9RISG1ꀿ��D�BPXWO���0 �zp$SK���2n DBT% TR�@' !^�Q0TC�� �`��DJ�4LAY_CAL�1iR� '��'PL	3&@�0ED`���'�Q�'�Q:�"d��!"�"1�PR� 
� �q��!#� T A$wq)$�љL@9$M?_3�Gp� %s?�4C�!&��?�4ENE�ax�1'�?_3!0RE�`�2�(H C�p o#$LC$$@3��B� K��VOa _9D6G�ROS�bcv�h�D��AMCRIGGEReFPAyS��ETURNcBo�M[R_o�TU�`)�2@EWM����G1N`��CBLA���E�Α�P��&$P�� 9�'�@�QU�C�D���0DO����-D�AS�3FGO_AWAYCBMO���Qm�� CSC0EVI>>@ ) HJ`1vsRBw���SPIhp�J�SP`wVI_B�Y��|S�UHSL�r*�XP$��avVTO3FB�\�dFE=A1v��SvTHS�+ 8Ɩ�DO?��cnpMC�%�d�P��)b�R����! `�,� $���J �c #fc ��faסߠebit�c�H�fa�"afWr��dNTV�fbV-pr��� ؃���g�s?�J�?�<�0��SAFE̕v�_SVq�EXCL�U�!����ONLd+�<sY�TktOT!!���HI_V5�PPLY_,�etw�]f�js_M8� $�VRFY_�#�O�� �v!1��s�b8Fc"�Q -�0� r~�_�:� �vGaSG� .�
$���@�A����U�REV�-�$��UN�0xK�vU��턍��@��l�i�!Xq����rEFf`I�2/��$FN�X$��OT�@jS$DUMMY
1ׄ1ׄ�����M�PNIG20C L����4���A`a��DAY�e`AD�iT� ��؃5��EF( $���1�0ѧ��Y�_3� _RTRQ�ݑ2 D_�Ot@R�Q:���'���Y� 21����~�jT|�8�s�¡3 0��ؑ �	�גS�U�@]��"CAB¡4��x��$��$ID��CPW��ӕH�g�ViW�V_Ӑ��0�DI�AG�q¡5� '$$V�@a�T�ǃ� ��� ��
0	�R�25���VE� J�SW������(���~����2ZP~�OH���P�P���IRs!	�B ��7�����Aᇀ��BAS9q�z ���HiV���4����Cנ��RQDW�MS�9���A�������L�IFE� ����10��N��
�ɵi���
�h��^Ui�Cm7Q�N�@Y����FLA�Tj�OV6նHE<���UPPO��w���� _6����vd�CT�6 `�pCACHE-�m���Es�B�SUFFIX�e`� ��@��R�؃6ԁi�qMS�W�7bKEYI7MAG�CTM%AH�x���A��INPU�}M�qOCVIEʠN�!8 m�� L�d<��c?� 	�q"��9��$HOST� !R�
0Z�0�Z�G�Z�R�Z�EMA�IL\ E�� SB-L��ULG2:"҃��COU��o�qT��0y�; $d��eSӐ4�IT1cBUFǂa�NTf Jj 5�B��mTC�dpA��s#��SAV<��҅�EK@b2W�Pp�m�PC�e�0ˤ��_0��"�`��OTRBu�
?P�pM�e���r��<Z͓DYN_�� E<��DtU� �U����TR_IF�nW�O��A�!=�0��/�Ӡ�#$@TCIKYD#&�L�A��p��K���/�DSP��6/�PC��IM<����sM�w�Uf�+�XE��p��IP�c/���D����TH0�|򲐙TLA��HS��A'BSCH���F��s�adk�$���oSCi��ʖ�1�!�!>bFU�I�DU��c��@PE���CD�	 ����W�R_NOAUT5O�!?��$����:�PS�C���C�"s�����ྥ @H *�L I ���jUs@�c >
1<1<G�<R��<��<79899P9��;E1R1_U1l1y1�1�1�1�2���GPR`�Hl2y2�U2�2�2�3��3E3R_3l3�y3�3�3�3ڭ4��� XTz�NaA <���� ��]V �jU��7���F�DRi�BT ��	���ò�17ò�REM��FQ̲O�VMb��5A�9TR�OV�9DTG�JMX#LIN�98PJf�'IND2@ʲ
^H* ^s�$DG
�X+��@M`ɵ��D��@R�IV�U̲GEAR�b�IO��K�2ʴN $��HY���_p�`�a̲Z_MCM��ñ�0v,�URwC ,��Wq?  �p?�0P��?0QE0op8QCa�aCOԐO`�D��n�P1av�RqI�QTz�UP2�p3E G���TD��os��S0�HQ�W�U����B;AC��F TP���T�Ł)]qG�U%��8� t IFI�� �XP]`+��UPT̢.�1MR2�5G���1�s�2LIxaFc�7��O�O�OF��ʵ�2_��N��_������M�F�O�MDGCL�F�DGDYxL	DHQ�D5Ѷ�Oɴ'c�E�H���i T��FS��F�I PแxqL`
�s�$E�X_wq�xwq1��E�Zwq3�{5�v�GsRA�P�4J ���tSW%�Ot�DE�BUG�#���GRt0���UZBKUe �O1  ΰPO`0��CԐ�t��MS�`OO��^�S�M�`EK����0_?E K ͠�P����TERM��L<��R��ORI`���M��ION�SM�_�P�҅�N������TAǉO����U}P�P� - �Ο2K$���L$�SEG�%pELT}O��$USED�NFI�<�Pt��� ��
�M$UFR��R��� 6�����`O�T��pT���0��N;ST��PATx����PTHJI� E0H�s� �=�AR��I�p��V��<�REL�r�SHFT =���nۘ_SH:�MO�"Ɔ р��5�O�a�0GOVR��r�&�I�j�dU� ^�AY��Q`��ID�MhS�� q� ERVDx�7  &�h2������!`ӥ��!`RCXQr�AScYM"�r�=�WJP�h1d@EhSב�����U'�������ђ�aP����V�OR���M@c��GRo��tQ ���U���l�����SѾE�R � h.�QTOC6�:�Q��OPbm���*t�v��1OA�RE��RT�r�O
�]⮒e�R��>����Te$PWR�@IM0ũ�R_���S��]� S�P$H|�U[�_ADDR�6Hr�G������vѷqR=p��8�T H�pS` ���#���#��_���lSEkq��S<� �sU $cP��_Dm0=���+�PR���PQHTT���UTH7�V (�� OBJECa!l(Q�Q$�6LE��)_�8�W�px7��GAB__A�Գ�S���I�DBGLV��K�RLp�HITE�B�GD�LO����TEM���%B�g�sSS�@7�HW��C���X��\�INwCPU�rVIS�� S���Di���j��j�~l �IOLN���Y} �@C�$�SL��$INP7UT_��$0���1P�@���SLp��aZ������IO@ЯF_AS]r[�P�$L�P���Q-�.Uƀ)�T��� ���z��HY�7T�-��U;OPZu\ `�r�6BBD�B@K���B�P 90�����K����&a�UJ�6] � v�PNEV�JOGk�n��DISBcJ7/нOF�$J8	7�W IT�'97_L�AB���) QA7PHI�`Q(mDypJ7J��0�p�_KEY�` c�Kk��0\s^ �@║V��{6�CTR<퓵FLAG�r;LGʴ_ �9`y8����sLG_SIZ��ԧPXp�FDI"Q�
 ��	��Xp����9����2@S�CH_H��R�� N�r`~����p�q��1�`UH�����L#�DAU%E�AP�k�ܴ3") GH�ݲz��BOO�Ra�t B3��ITp�3g$�`/�REC|*�SCRN� /�DI2.�Sl�=pRGMb�0��,��'����"���S����W�$�$'�J{GM7MNCHF��'�FN�6K;7PRG99UFG8W�G8�FWDG8HL~9STPG:VG8`G8n G8RS�9Ho�c;$�CY��3&�'��p�'IUG�[4�'H��&� <�2N2G+9�PPORG�:0�%�3P/6OC$�J8�EX#�TUI95Ii�#�B�#�C3�C 70;11���AC�'1�v�!NO�FANA�6��`VAIQ ��C�L�a��DCS_H!I	�NR��MROSX�a&VTSIxWjXSvX�(IGN"��481� � `UUDEV$��B�U`��b� _�T6�B$EM�[ᨽk�3A��c� @_���e�W�Q`m@19e�29e39ae}Q��d ����{�5���%��IDopX�.�4�=aX�&���fSTs�R4 �Y�p1��` c$E�fC�k��F��fp�f\тD��e LL� B��pW�)�� �C�����PЄ��"�#_ f ���V����!�s|�C�g ����CLDPs���TRQLIi � �y�tFLG�b�p�a�sb=QD��w=�LD�u�t�uORG �2�r ���8��ç�ҙt0�h � 	�u�5�tJ�uS��T�p� s��!�����RCLMC��<�N�������`sMIН�i d��yaRQ� s�DS3TB���` ��!�'�AX��� *�C�E�XCES�� ��MO���j�P���k���Nџ�k���_�A���A�S��pK�ʴl \L��$�MB>�LIw��REQUIRˢ
��=O�DEBU`B��LSpM�m��4�Z�h�������ND	!�ǰ��n�����DC�B$INeЫ!$�� ���PN�b�C��PST�� on��LOC|fRI&�|eEX�A��}a�^��ODAQ�p
��$ON�RMF �@`��iRrJ@\u�����SUP��R!F�X�IGGz! q �s�Rs���Rs4FRtR��%�cι�s�޸s��ΐ<�DASTAg*�Eq�E�t�T�N�Rr tN�+MDK�Ix�)YƎPd��a�H/�"dĸ�<Ue�ANSW�!d�(a�Ad�D&�);���ܔ���s ��CU�"V���p7�RR2���t���Z���A��� d$CALII ��GAQ
�2���RINP0�<$R��SW0ʄH�y�A�BC_�D_J2SqE4��X�_J3s�
m�1SP?�< �	PmԔ�3����������Jy��Մ�V_�O�QIMy���CS�KP�z��:S�J<!��Q�3��3�)�$�_AZ����e�EqL�Q���NTE��"bu����7���%p_N��v����a��4�䛒w��DI{����DHc�����x� c$Vв��a$;1$ZbN`b������yH ��$S v�TqACC�EL�QU�ׁd�I�RC��T?�T<�a�c$PSc��rL������s��z�x�BP{�PATHZ����p���3���f�_@6a$� ��M`C���k�_MG�!$D�D${�"$FW���=�`�@p�k�5D}E^PPABN��ROTSPEE�:a��p)�:aDEF�!�k�$USE)_�SP��CO@S�Y� 6� ��YN� �A� ���{��M�OU!NGO� O9L��INC��,��]D'�=��(�ENCS�#����k�%���IN�bI��>����)�VE"Ӡ2�3_U�b�LOWL�QI@���pi�D,@�����Wpir��C���MOS�P�ӔMOܰ����PE�RCH  �OV � �1'|a<#�a��� �a2�m"�,����P��A��%LT��З��ך����&�TR�KE$�bAYLOA ���"�� 1��53-��`S�RTI��K�`MOM�B'���2����\
�3��9b5��DU����S_BC?KLSH_C��5 &D ��°4d�:<+�CLAL`�p��A0���5CHK�p:�eSRTY�@(� �@�e$�<�_�c$'_UM��=ICJC$�SCLWD� LMT��_L6���pE��|GEvM�@�Ku@���E����Ц1
� �Du(PC�B!u(H��;�(@EC̺�]rXTk�6CNE_%�N�S7V׃S�P� g(V��c|V�Qȟ�{UXC!`HMSH �c%�6l$�{1{�`2���U��$PAGD&;_PFE*3_�pd@�6% �q3)dEJG0xpy�c�OG*Wn2TORQU� ��#� 9l ��"o1l �b_	WY5 4_�e�eT�eI�kI�kI�FE��a��x]�. VECZ�0!���"r1(~pu�<2�/uJRK(|�mr`v��DBL_S�M7��M��_DL�GRV�d�t��t�qH_�S�s����zCOS�{/0�xLNop
�+u����@��aH�6��a�uZ��&�qMY����rT�H�}��THET0�NK23�т��CBֆCB�C  �h����d	��	�ֆ�SB�'��GTS���C��,��S&��P�S�6�`�E�$DU @И��
�G������rđQ�2�$NE䂗�I�(C�2R���$��ŁAɅ����u�x�qLPH�uВ�ВS'�C�6�C�E�ВT�Pm�W�t���V�V	�T�,�V;�VH�VV�UVd�Vr�V��V��H�-�3�+��QJ�H�UHV�Hd�Hr�H��UH��O�O�O���*�O;�OH�OV�O�d�Or�O��Ot�F�В��R�6�W��SPBALANCE�Զ�ALE>�H_ɅS�P��'���6���E�PFULC���½����E���1uLUTOy_@=eT1T2�V�2N�1q�)�6���@:1�������U1T� �O{�c�`INSE9Gq��REV��ΓDIF�%��1vl����1w� OB���1�sg72x`)�A�t?LCHWAR���AB�Qi5$ME�CH�����(FAX1P�D,����Їx 
-�aO�|ROB% CR�"o�!R=��MSK_��9�_z P !�_� ARV����$1zR������4����I�N|��MTCO�M_Cp=�{ �  ��v$N'ORE�������o| 4�`GR�b��FLA|�$XYZ_DA�B`��/DEBU?� ���$�} ��$�COD�1 o�>2��90$BUFI�NDX� ���M{OR��~ H�� W0e��6��5�4�ҎJ�&Q��@TMA���g2G��� � $SIMUL'`v�X#��#OBJE��A�DJUS1$ AY�_I>az(DROU�TG`>�W0_FI=��T�`�	� �I��Ф`� ��в�:�%D� FRI�3�MT�5ROg`�E�a>� �OPWOnp����,|�SYSByU⠙�$SOPȇ��1U��PR�UN��<PA��D;�s _m �B1���ABc��@m IMKAG�1�ฐP��3IM��IN�pd~�RGOVRD�- oPq�xP�ЃL_	ЄQ�<BWPR�BXP���AMC_SED��� �@N��M"�A�0MY19��A��SL������ x $OVS�L[�SDI� DEAX@SR&OS�!p"V�`m%Nw!�aj� u#�'�(%"	�U2"_SE9T�`��� @�`�"L6�1RI�0
�&!_��'�!�!g���\/ lP ���T��<`ATUS~0$�TRC��� ��/3B�TM87"1IY#$4p�A3 ��� D��!EmV",2�E��-1p�� �0-1EXE30@)A!�2�2f4�#�� ̟�20UPI�1$�ИXNNX7q#$�q[9 �PG��� � $SUB�!16��!!1�#JMP�WAI�PPz#9EL�Oy@9��$R�CVFAIL_C��RP<AR�  �)�Q�jPATs��E��R_P=L�#DBTB<anR�RPBWD~F�UMl`�DIGT�<���@DEFSPH� �� L��3��@_8�@7�CUNIr]7��@�1R�0Ҥp_L���P+1��
@���� k�e`�q� J���N��KET@R�`W��HPP�B�� h~B ARSIZEw��:� I�QS/ OR~�#FORMAT���DCO5 �Q~�EM2%��T#SUX� �"��BLI�B�� � $��P_SWiI�ЏA��AX�@��@AL_ � �$�A���B!��C���DY$E�1��,`C_�A� �� �@�d��(aJ�3r����TIA4�i5�i6��MOM���c�c�c�c�c��BP@AD�c�f�c�f�cPU
�NR�du�c�u�bER a�� C$PIǖoe�� od�tWu�sWu�sWu���vm{ �r�[!P�j!�{�$�6�SPEED��Gb�tQE�D�v �DQE�@� �v��x�A8��AQESAM����pZ��w[�QEMOV�� �����Л��������@	1�䶄2��� ��`Ƞ�%`�H<Т�IN �%`>�����QB��2�	�2�R�GAMM�~Ʒ�I�$GETH���;D_d��
1�OLIBR�1GrIT�$HI�0_�;0��ǖE��ԘAΞ��LWɝ���3��\[b%�MTN+aC�E�����  $�PDCK�$�;_ =�� ��$bph$a؅���c���f��)c W�$I� R"�D��0���1rD��LE�����!�[h�n`MS�WFLY��T�И���Pq�UR_SC�R�3`�-�#S_SAVE_D�~��3NO_`C�!�2`d~� ��ojXv��qy��0� �ۻN���v�̀Ja ` <����љ������� �x�v��|�x�6�Л��11�PM2u� 7� ��YLQs�� ؇Pу�ɣ�Ǟc��B��W��w����Ґp�����M��(�CL'�(aC&"l�"&�qΉ�PLMo��� ό $���$W~���NG�ya~� 8d|�?d|�Fd|�Md�@@��᪐c�%`X9P	OGc$aZ��P@ ��G� pB ��ʣUv���ҿ�����_a_�� |B oi~��i ��c��c~��j���患jE@ ���U��U���\�z`��P�Q�P�M� QU_� �{ 8TPQCOU̡n^ QTH��HO��nc�HYS�PES��Fb�UEN�t��POd�   ���"sUN40*� 
@9O���� P����oE`�}3GrROGR)AG1��2�4O����xR���INFO�ᇗ ���� ���u��I#� (R�SLEQ�vK�uK H�����D>@��Т�O�����sƑE��NU��AUT<���COPY���0(�j!��M�N� ��m�C� �QRGA+DJ�ᚓRX�RC$9P.�.W,�P,$�.�s�#E�X�@YC���AR�GNSD� � $ALGOz����NYQ_FREQ��W=��v��T�#LA��ѫc=��u�CRE�0�#� IFl�#��NAc�%��_G�&3(%���E�LE-@ �jbE�NAB�ҡPEASI_!|���N"�q���&cBՀ��I ���`�qf�_`��"AB�!�K`E���pV��'BASUb�%�����0���0$�!6��� X �" 2� ����@>62=7;QX�ޠR5Pi6�B�-PF��ROGRID�13CB�P��wTY`#�OTO����@��_$!HZ�2C$O ����9��[@PORqC�3\Cv�2SRV )	D6FDI�PT_�p#@�5D��?G3=I"P?G5*=I6=I7=I8!A�A�F������$VALU�#q�r$BR�A>��| [%������3!n��PAN�p�vS0 R�0�Qn�TaOeP`���$SPW��I�1:TREGEN8ZMROcX7�s�v���FI�TR�#1B8Q_!St��WMP�#Vѵq�U�q<!GRTb�Q��Slì� SV_HƩ0DAY�P�PS_�Y�����So�AR�Y�2�+0CONFIG_SE_�PB�n�d2���G�5� 4�W�?�vv[�6�PS�~��� @W�MC�_Fl�|�a�L�~��SM����a��bNs����c� �,R�FL�Г���Y�N�`|Mf0C���Z9PU��LY�ᦛ�ODELA4pb�Y���ADY� �QSwKIP�ŧ ľ���O��NT��o1^pP_����}w`��ҵ� �w�Q�y�Q�yV@�zc@ �zp@�z}@�z�@�z�@z�z9�q�J2Rf�Z��fbEX��T� C�n�C��0rC����q�0RDC֩ ���R塘�M�ͅ�����f�w�RGEA �R� ]��E�D��ڝ��ER�a^�C~U�M_C�p�J2TH�2N��4� 1�[ t�EFI�1��� l(�4�\#��Υ�TPE���DO �]�����T���O3�S���Ւ��~��&�2.��4�F�X�j�|���
��3.����ß՟�(�����4.��.�@��R�d�v�����5.�������ϯ�����6.��(�:�L�^�p���
��7.������ɿۿ(�����8.��"�4��F�X�j�|Ϡ�SMSK��#�
�'�bP<D��1REMO& ��f`�6�V4�IIOT�I���PI1��POWER�� �6�pa����S ���e��$DSB � �!T/pC��B^t�S232:ն� �*�DEVICE�U�". t�RPAR�ITY�.!OPBI�TSFLOW0`T�R�� R+P���RCU���r UXTAS�K�RINx�FACp��1"��0�SCH����b�`_sC�����POM�tbPGET_�@�b� g0��m�P[���� }!��$USAp �1���� O�`� p��'`���_ON�qP����WRK�����D�P���FRI�END 1x $U�F��#w�TOOL�~�MYH�`t�LENGTH_VT��FIRM`���U E|�е�UFINVw �RGI�MAITI�r��X�zq�� G2 �G1@�1U���+�0_y�|O_�Х���#0� ����@TCs��D� �G߀1#b`��`�����bo
�0.%�S0#�R �����>��X ��v0L�T�H�0���&����)$W�0��EDRpLOCK�6'Aqwp�QUi�Q	$�20���4�.�:��1F�5�28�2�38�3F���G��! �����S���SV�P��VVV@�`b`���b��so:�|+e p�qP]P�! @��S��U����A9@��'PR�P�&��SS��q� �q���2� 0��0�20�haV#�������E U�{r
��S^��� �c!RA,Q{2$P`N��`�BHAn�L��rw2/THIC.� pap�C��TFEREN�1t5I�@H.�w1I08��3��K0G1�(�4����9�r��6_JMFGPR�`}q�b��C� <q� *R �}r�C �-F{� ���ҢA  2� ��Sx����	d' �$��Du��Ep�C$Pn4�CDSP�F�JOG�P�p`_P�q:�O�1Fu��� L�7KEP��IR�A�D2]`MUAP&�!E�%P�4�S`�@��R�PG:VBRK�`�5�0n0I�� A aR�clR�Br A�R<�C�@BSOC�FJ�uN�UD#`Y15�q�$SVDE_�OP9dFSPD_WOVR�a<pC�`L�R�COR�W��N��b�VF�1�V�@OV�ECSFjP`c�F3f��!�CHKh��"LC�H2rFuRECOV(�T���@W"pM�P�eF�@RO8�Q�@_h0�a0 @���VE�R�p��OFS��CN@��WD�Q�d�Q�QX��U�PTR,� Ѿ#@E_FDOVMOB_CMb�	pB�@�BLs"�B+rs!�$V@�	��� ucbG,w?XAM=SpZ mu�b�_MCpE�ހOӹ`OT$CA�@ހDhR�pHBK��6�q�IO8��upсPPA�z��y��u�u�pҹbDVC_DB ��C��1��D��b�![�1c��s[�3c��`ă�U��@�QUK�@O�CAB�@7��� �ch� fx
�OzpUX�6?SUBCPUr2�@SQ��sUt��*#��3#Ut���Q$HW�_C��D@pH�A�.c0�$UNIT�uTo�h�ATTR�I-P|��@CYCL�ycNECA��SF�LTR_2_FI`�4�خ����1LP�K��0�0_SCTvF�_h�F_r�����FqS��Mrm�CHAQ���<�Lr:�;�RSD��`�҅Q�3s1p�_T�jxPRO��s0�E%M��_�`iST)�:!� )�C!��DI����4RAILAC4Q��Mz@LO�P���T7t� ���!���s+PRE�S�10��C7���	�cFUN9C�R�"RIN� s�02�Ġ:�/�RAK��� �pc�p�tc�W3AR�3�pBL|y��A��������DA`sPd�θ����LD�� �P���o1m��!��aTw� �vcc0$��gRIA���AF�P�Aä`GŶ[�S�ʓMOIs�vD�F_��Jc��C@LM�OsFA��HRDY.�ORG��H]�v�2�ְ��MULSEP��-S�L!��J�Z�J�Rg	kFAN_�ALMLV,��W{RN�HARD`����� ��n�2$SHADOW`�0���AMU_�`�6AU�� R.�F�TO_SBR9��յ@��h�9�|B���MPINFa0!~������g��p��`|A�  d�m$!�$�� xB|bA}@�� �2S�EG� �C�P%�AR�@���U201躰?UwAXE�GROB�F�W��fQ_t�SSY�rP_�hP��S��WR�I��8�*!G�ST�R�E��gP�PEj�HK@A�oҽ B���a���!�P�pOTOr��K@�`ARYn3`+�䡘�UA�AFIHP~�C$LINK���~1K�/!_��at@��!r�XYZ:�:}�5��OFF�`J�)r�f�/�B�@/�����a��3���FI@����:1�R�T/��D_J�AIB�RW�e�0���S�TB!��2YC��.VDU�b?�.��TUR�XÒ�9��X���pAFL�0 g`ǃ2� ����8��R�a 1�K@K�@M�4?�9����"��cORQ���Ai���3H� EP�0���!�`-S�ATrOVE|�2M��1�Ӗ�� ��IГO��j� �E4��H��1}�@ �d��1�}�%�Ә%��AER�Am�	B��E��1@�]$A!c0��[���7�ձ҆ձAX�cIBձ��Q� L�%���)���)���* ���*�P�*���*� �*�*1H��&���)\0 �)\0�)\0�)\0�)\0 9\09\0/9\0?9\1�P9DEBU@�$�;�Gӯ� A�bn�AB�է�q�Qv[@Ġ�r
 Bl�7!CEb�OG�OG ��OG��OG�QOG��OG �OGM�^ G����LAB��A<�I�GGRO��A@��pB_��D&���S�����F,QB(U��4VAND� ��R$��w�U!��qW �q��v�XƱ�XL��v�NT'���ПSERVE�P��� $��g�Axa!�PPO�b��p%��Q��S_MRA�� �d ԰T�`xdEcRREsC�TY.����I�pV��#2aTOQ�$�Lc�$���Eeh�SW�� �� px ,P�d��_VA1^2�!�d���d2�k!2�f�QW�� �@@�Q��s$W���fkeV����$���w��dd�SOCƱ�� � kCOUN�T�� �QHEL�L_CFG��� 5 B_BA�ScRSR AB��#�i�Sj��cpU1�U%bq2�z3�zU4�z5�z6�z7�z98�wVqROO���p�ݐu�NL��dAB��S͠dpACK,FINpT�4��e���.��_PUՓC��OU�SP��guܡDr��v��чTPFWD�_KAR7ac aR�E�T��PG�ܱ��QUEm���}���A�c�I�/CCss�ڣ?�8v�at�SEMR�	��b���<�.PTY%�SO�!DDI1����C8с�'u�_TM�P"�'NRQb�s�Eߐ C�$KEYSWI�TCHڣ��D�ڄH=E��BEAT�����E5�LE6b����U҈�F����SI�DO�_HOME�OO�REF]PR��"����2�CԐO��`qa�O�P3@�&�IOCqM_�YA�Av;HK�� Dp�o�ORESUbςM��x��ooFORCs�nʳ @wOM6� � @
D=Â�U��P4�1֦�4��3֦4���NPXw_ASKr� 0qp�ADD{�Z�$S{IZa$VA2P\�u��TIP��
۠A���``_��H���]�S�C�C2`�y�FRIF��pS0��˩�i�NFe�
��dp�� xx SI�ObTE�P�SG%LѱTY� &���x�C��ҰSTMT�2�P!���BW}Ӵ�SHOWř��S�V����� �	aA00vTT�ߠ\�@�\��\���\�5Z�U6Z�7Z�8Z�9Z�AZ�W�\�ʠ\��A]ƀ��\���_�O0�f�1�s�1��1��1��1���1��1��1��1���1��1��1�1�1�G���f����� �ɉ��ؚ�Q �ش�� T����2��2��2��2�2�2�V��f�3s�3��3��3���3��3��3��3���3��3��3��3��3�3�4��4�f�4s�4��4��4���4��4��4��4���4��4��4��4��4�4�5��5�f�5s�5��5��5���5��5��5��5���5��5��5��5��5�5�6��6�f�6s�6��6��6���6��6��6��6���6��6��6��6��6�6�7��7�f�7s�7��7��7���7��7��7��7���7��7��7�7��7�7ԃ��A�P��UPDJ��� �`� {r�aYS�LOKr� �  #�i�f����S �4R@U5;���p�R@8F�!ID_L,e�h5HIc:I���P�LE_b��4�$�	��&SA�b� h�`�0E_BLCK��2���8D_CPU�9$��9�c3�?�4x�"P]�R �|`g
PWp�q FALA��S�aKC\AUDRUN�ErAJDrAUD����E�AJD�AUD ��TBC�CJ���X -$�ALE�N��D��@?�RA���R� W$PI��F)1�A�42WMp]�h�C��.�ID� jQ�&\TOR�@>[Dx�a0S��LACEB��0R�@c0R6`_MA�	�MV�U]W�QTCV�\�Q]WTn��Z�U�Z@СKT�a�U]S�aJA�&
t$Mdg�J��D�RLU9a]U�A2A�`<��`RaKS"PJKefCVK�wa�wa3ic�J0�d{cJJ�cJJ�cAAL{c�`�c��`�f4�e5�B�QNA1�\�`�[�P.TL'P�_��>��!�@Is�{ `�0GROUN0��g�B��NFLI�Ca�=pREQUI;RE
�EBUJ��AfY��P2�X��@]vx�A�G�� \m�/APPRipCT��P�
��EN�xCLO��yS_M����y�LU
�AL�� �7�MC�R�P�B�_MG���CF��0$��␉P%�BRK#�N�OLS�%�2�Rc�_CLI%�i�S��Jr�e�P�diP�ciP�ciP�ciP�ciP6��߱���8B����A�t��# fr�B�A ��A�PATH
�#���#��H�N�xp�`CN�CAt�i��r�IN�BUC-P1y�-C�PUM��YPl���l1E�@���@���`~o�PAYLOAa��J2L� R_ANx��LG@��ߙ���$�R_F2LSHR��%�LO�x�)����7���ACRL_@�v�i�r�ה�BHA0ζR$H$���FL�EX�s�AJ�E� :�O�F]Pȧ�ߤ�O�A]P�O�O\F1ߡ-�A�_)_;_M___q_q�E{_�_�_�_ �_�_�_�_oH�e�g $cedU�w�,o>oPoޡWjT��F�Xl�bce ����ne��zo�o�o �`�e�e�e�e�o�o�o�y�J!t� � �-?Q��� AT�Z�eq`ELȰ �*�lxJS��spJE�P�CTRr�U�TN�v�F(�]wHAND_VB���M0�7� $��F2$��s�b�<2SW�ӴA�v�?� $$M��R>���O������厂�Ao0ܐ�n1$��QA.�10@�AN�A]�P/�/��0@�DN�D]�eP=�G]@��STB�h��O���N`�DYt@ �p$��7��}��ߡ �:�ޗeg�����d�P������Å̅Յޅ8��Ӓu� �ത���"��q�!ASYIMM��fpM��`8h�:�m�_SHrw� ��{��蛟����џ�Jꜛ������.g�_VI����s>	 V_UNI/�$?�'�Jfe6"d6":� :$Q�G$k&Z�`m����|����%���������@�pHH@�r�̙��!EN��
�DI�]���O4�� !sS� O�>�I!A���Q�819@�3F3�08�O��:B�1� � ��ME����a2�"HT� PTq��8��1pt�p��8�1�9T�q $�DUMMY1G�o$PS_X�RF�ֽ�$�6!ALA�#pYP���2�3$GLB_T��5E��01�@��Y�'1� �X�p]w�ST���spSBRM�M21�_VbT$SV_�ER�OWp_CwCC)L3@_BAɰO;2� �GL  EW$q� �4+p�1$Y�ZB�W�C[`$���Ab0҂�a큤AU�E� ���N�@v0E$G�Ii�}$�A p�@�C�@$q� L+p��Fr}$FrWNWEAR��N_�FLY^��TANC_�@��JOG?��� ����$JOINTx�!q��EMSET$q��  �I3Tʱ��SpM�U��$q�����MOU��?�spL?OCK_FO9����0BGLV\�GL��XTEST_XM��p�QEMP�P��xb1B�P$US~1��@� 2�sp�C@a��b���P@a�aACE�pSa` $KAR��M3TPDRA8�@~duQVEC�f�yPIU@a�EaHE��PTOOL!��cVv �RE�`IS3�r�d6ÁU�ACH�P�S���aO[��3�42��PSI�r � @$RAIL_�BOXE�!spR�OBOd?�aAHOWWAR��0q�0�aROLM�2Vu�р�dgr��p�T�a���_�DOU�R� H R^cI2���P_$PIPfN�� �br�ag�@a�q�B��}OH0 � D�pGLOBA�6��P����3@�r8�SYS�ADR7�� �0�TCH�� � M,��EN�"1A�Q�_�Dp���3� V�WVAd1� �� �`�B5PRE�V_RTq$E�DIT��VSHW�R��KFԀ���A��Ds0
���HECAD�� �����KE�A�0CPSP]D�JMP_�L 5���R��#4���e�I`S7�C}�N�E�`8�s�TICK�!�+M5�F�HNAA� @�pc��Վ$�_GP��v&@S3TYj��aLO3A���F������ t 
���Gv�%$���D=:K@S�!$,!� �x1E50FP��S�QUx`�B�TEsRC�0��TS��� �&AW@�ר��׈x��aT�O�0�3c�I�ZD�AE�1PR�OC�2Ѣ1�pPU�#!�_DOQRo�XuS�PK 6AXI �zsEaUR�ɳ8� 7p��.����_�`@��ETA�P�R�����F�
t�R���l ����� ���榹���� � ��0�ڵR�ڵb�ڵr� �͟��*��
��s��C)�k}�����SSC@ � h�@DS��a�03SP20�AT`���⡠�o��2ADD�RES�cB��SH�IF��7`_2CH�7�*�I:@X��T�XSCREE��z���TINA�CPk��D��B��C@� TU�z@Ţ8�yA�V@���7���Լ�RRO; fP7����W4v1UE$4� �� �Y��0S�A8�RSM<���UNEXk� 6"�� S_�CB�%2�E�`�%B�C�R��o 1�t�UE{���,2�B��ѠGMTJ~ L�!�f@O�V��$$CLA<� ������0|����VIRTU� �����ABS����1� �� < �� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/??�+?=?O?^;���AX�L�����+�  �p4INy?�1o4��/_EXE�8�0�6_UP�м1#����LARM"�OV ���2l4LM_�P���d^?BOTOfOxO��J0O�O�O�O�O�M�, 
6�_j6NG�TOL  #�	? A   L_^[��PPLIC��?���0�P�Handlin�gTool �U �
V8.10P�/11  S-�C�(
yaSW��R�����
�QG
F0�Q�U�᪚п
1232�T���
`��
X�{s�Z�s`~��7DC1�P�\�SNone  �EL@TFR=A_ 4�YWbql�PpQ��TIV�5t�S�3�cUTO��� A�4�9P1�GA�PON��n��`O�UPL�p1I� �`&g9�`]UB� 1K ��
0x0|0|����s��1�s��� g��UvtH_u�r�zHTTHKY���cu��� �#�}�G�Y�k����� ����ŏ׏����� y�C�U�g��������� ��ӟ���	��u�?� Q�c�����������ϯ ����q�;�M�_� }���������˿ݿ� ��m�7�I�[�y�� �ϣϵ���������� i�3�E�W�u�{ߍߟ� �����������e�/� A�S�q�w����� �������a�+�=�O� m�s������������� ��]'9Kio �������� Y#5Gek�|Bu�TO6P�o�cDO_CLEAN�o@t#_NM  ;[_�Q/c/u/�/�/4_D?SPDRYR/?uHI�`/-@@/?? +?=?O?a?s?�?�?�?p�?�?�?<xMAXrP ����g�1X��Q��b�Q�bPLUGGp�`��c�ePRC� B- �+�/�?WB�O\B�/@tSEGF�`K�O�G�A-/?/_�_+_=_O_�O�ALAP�/�N�s�_�_�_�_ �_�_o!o3oEoWoio|{o�cTOTALF|HI�cUSENU�@��k ��o�BpR�G_STRING� 1�k
�kM�`S}j
q�_ITEM1v  n}m6HZl~ ��������� �2�D�V�h�z����I/O SIG�NALuTr�yout Mod�euInp̀S�imulated�qOutތ�OVERR�  =� 100rIn� cycl҅q�Prog Abo�r�qȄSta�tuss	Hea�rtbeatwMH Faul\�e�Alero����� ����ß՟�����/� �{�( 2���������ȯگ� ���"�4�F�X�j�|��������ĿF�WOR �@{��p�ֿ$�6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h�z�PO{P���� ������������/� A�S�e�w����������������DEV��D��1�k�}��� ������������ 1CUgy���>�PALT\�� ��"4FXj |��������//0/B/T/�GRI@{�! f/�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�?�?z/�`R\�0A�/
O XOjO|O�O�O�O�O�O �O�O__0_B_T_f_�x_�_�_OPREG ��PHO�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@����$ARG_��D ?	����q��  �	$��	[��x]�w����yvpS�BN_CONFIOG �{ցՂ��qCII_SA_VE  ���q��rvpTCELLSETUP �z�%  OME_I�O����%MOV�_H9�L�R�REP�3L��pvUTOBA�CK$��}�FRA:\�[c ���V�'`;���W�� �� �x�]>�P�}�pt�����愈���� ����)�;��UΟ g�y���������L�� ��	��-�?�Q�ܯu� ��������ϿZ�����)�;�M�_�>A�� dωϛϭϿ����ϲ��INI�  ��u~��MESSAG�����p�ODE_!D>��͆9�OF�H�޶�PAUS��!�~�{ ((O�r �߲ۜ���������� �*�,�>�t�b�������{ԅ�TSK � ����Ϲ�UP3DT?��d5�U��XSCRDCFG� 1�v������|��� �����������e� 0BTfx��� ������|rs��GROUN)�|i�UUP_NAf���{	��R_E�D�1
L�� 
� �%-BCKEDT-Cz���[��t]�-����Z��r��W��r/  ��_%2h/y�F/�/<"��t%�/�/C/U/�/y/a#34?�/�? �/�.]?�??!?�?E?a#4 Op?MO�?�.)O@�O�?�?�OOa#5�O <O_`O�.�O`_�O�OO_�Oa#6�__�_,_ �.�_,os_�_o�_a#7do�_�o�_�.�o�o ?oQo�ouoa#80�}h�-Y��Aa#9�lI�4��-%�������a!CRg/�o�&��m �Z�����I�׏U�?NO_DELas�GE_UNUSE�_qLAL_OU�T ��>#tW?D_ABOR���T�ITR_RT�N׀l�NON�S��.�1�CE�_RIA_I)�j5�y�FF����.��_PARAMGP 1����?
���.��Cp  O���Q��Q��Q��Q���Q��Q��Q��Q�ҪQ��Q��Q��Q��7  D DI�p�����y�ͅ�둴�� D��Ѱ���"Ѱ*��1Ѱ9���@�.?�y�H}E��ONFIG#����G_PRI 1���Ё$��S�e��wωϛϭϿ���CH�K��1�5� ,5���%�7�I�[� m�ߑߣߵ�������@���!�3�E���OF���찫tCO_M�ORGRP 2�֬ h����� 	 �����������누�̣������q? ����p�`�;Kh�:��Pa��!��a�-��������.
��
��r�q@����.�`M/CPDBc��$�  )cpmi�dbgN�� �:_�  /� ��p������O  �商�4-���+��v�����gHf���f��/��/� mc:�,/T/kDEF �"(�)@ c�ebuf.txtp`/�a/}�_MC��mu ԰ d�%�#���-���!5�Cz  BH�B����B�pB���6C�B?�r-C@�F��C��kCw*��C�"�D@O�C�0TDK�#�Z=E4�E��D�l�E��dE/BE��C	��)4���C<	k���~k��������A�x��g1\Q�DD�i�D@Z=DN@ �DE�D�  F��E�oF`[/R�> �JBEL@�Gb��FO�\�G�L��:�  �>�33 ����;  n��;�#5Y�E��; Aa��=L��<#�
�E�O/�"RS�MOFST �.���)T1��DE� �� ��
,�Aj�;��B�O�O^�.TESTy"._�v�R��g��_%6C�4�@���� A��A62��;0Bl�;0C�(@@c��j�:d[�
�QI_���]��QT��FPROG %,���o�UT_IܑZ@䖏��d�KEY_TBL � 6��
A� �	
��� !"#$�%&'()*+,�-./01234�56789:;<=>?@ABCy �GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~����������������������������������������������������������������������������q���������������������������������������������������������������z`L�|��kp�z`ݐSTA�"��T_AUT��O�e��V>�INDTO_ENB+���ROQI�;�T2��t�a�n�v��XCˣ 2�j���8
SONY? XC-56�_	B}�u��@��Ͷ4( А��HR50
���+�y7=�O�Aff[��o��ß �����՟ �0��T�f�A������w���ү�����f,T{RL|`LETE��� w�T_SCR�EEN ,�_kcsc��U���MMENU 1u <*�o�� �����Sǿ�&� ���\�3�Eϒ�i�{� ���ϱ��������F� �/�Uߎ�e�w��ߛ� ��������	�B��+� x�O�a������� ����,���b�9�K� q������������� ����%^5G�k }������ H1~Ug�� �����2/	//�A/z/Q/c/�/�)k�_?MANUALÏF��DBCOe�RIG�4�5�DBNUML+IM��s`d�UY`�DBPXWORK 1 fk�_[?m?�?�?�?�]DBTB�_)� !�_�Q��PK4�!_AWAYz�#:�GCP �R9=|P�6_AL0-���2�"Y6��P�(_�DBG 1"ZY�I�,�K?�O�SrO�O��8_Md�I)PL@|+`�CONTIM3����T��F?I
��eTCMOTNEN�D�oSDRECOR�D 1(fk �<�O�SG�O�Qm_ �[B�_�_�_�_xX�_ o_4o�_Xojo|oo )o�o!o�oEo�o 0�oT�ox�o�� ��A�e��>� P�b�t�������+� �������:���E� ͏��������'�ܟK� ՟o�$�6�H�Z�ɟ~��i�w����@37  � $2201		! US�@ܯ� ��o�$������ es�erved fo?r SETUP��������ȿ7���[� �TN Menus� %ASM #2 ��4�Fϵ�j�U�c�����@OUP) $w040�� #3�� ����Y�����D��@7��$Fc�E�|ߎ�����JTOLERE�NC DB�IB@L���� CSS_D�EVICE 1)>�9  �6� �)�;�M�_�q�������C��LS 1*���������!�3��E�W�����PARA/M +`Ii�����_CFG ,�`Ki�dMC:�\��L%04d.'CSVh�H@c��i�YA"�CH zH@��Oi�Q���'��2�!~l@0�J�PѦ�RC_OU/T -�;m@k�~��SGN .�5�?R?114-M�AR-22 14�:45"���? Tnu�-)�i�*��\�o���Im��P�u�G�=��VERS�ION �
V3.1.0�L�EFLOGIC {1/�; 	�(�@0����PR?OG_ENB!OFRF�UL١�%�6��_ACC6(A��.C�7#WRST�JN�@�&��MOp,(A0E{!INI� �0�:�5?1 v&O�PT_SL ?	��&�"
 	Rg575i�� 74�)�6�(7�'5�21�82�$�6?��$TO  �-@�?�]V� DEXd'd?U��3PATH A�
A\�?�?O��KIAG_GRPw 25��� ��	 E�  Fw,D FAD�`QC��@IC@��nOLkA��ЗO�NCeE�Cl^OCkI$�C��C� �B�m�If�362 6789?012345�B�'�  �cPA����A�=qA��A�33A��z�A��A���RA���A��P���JPj!@�\@p	 GQ��A�2����"�B4L�ѨD�(j!
R�P�{A�P�P���P�P�G�A���\A��A�Q�*?_Q_cT�*��T�)�^�PϸP�P�� P��P��P���A�ffA�P�#P�_�_�_�_o�X_�PZ@`U�PO�
�AJPDP>$P8
P2@`,�lWoio{o|�o�]`��A[�P�V�PPPK
=A�E�A?P8�w�A2�P+�
�o��o�o�X��`��$PLpxPqPj�$Pc P\Q�ATPL��bt�� ��TC@R�Q3a�aKq��p^M=�G�z�>�8Q솅^M8��=b��7�Ŭ��^M�@ʏ\ʆ�p�4օE@[PAh	 ��C@<�C�<�t��=�P=�h�s=���~�C@;7��
.�<#8�[� �?+ƨC�  <(�U�w 4Ƃ���r�����~���@
"? fE6���8������9� k��0�ʟ@�f�H���<��~�?Tzᾦ;�dʥ^M�{��G�^N cQ����^Nx��7���C��O
�@�CkJ=C��CCk�^M�����|����`K�
�׿M�ED  Ew�� ��D+�	��C��O7�j!8���6з��3��V�?6г��G7�����İR��=yġ�C&=A�����#Ϡ����{������I ACT__CONFI��6������eg�� ASTBF_TTSd'
)B�C#t��U���MAU^ \/��MSW��7���_P��OCVIEW�i�8��	 �� �����*�<�N�I ��~��������g� ��� �2�D�V���z� ������������u�
 .@Rd���� ����q* <N`r��� ���/&/8/J/X\/n/��RC��9�5v�!
/|.�/�/�/�/��/#??G?[�SBL�_FAULT �:�*��a1GPMS�K�7t7�0T"A �;ٵ���M�C: �C�O�:|#P ��OO1OCOUOgOyO �O�O�O�O�O�O�O	_8_-_L� ����1ORECP�?�:
�3 �_���?�_�_�_�_o o,o>oPoboto�o�o��o�o�o�o�oI_��U�MP_OPTIO1NK�m>qTR��L�:q9;uPMEJ�.�Y_TEM�ï��3BK��p��ytUNI��MՏq���YN_BRK �<��y8EMGDI_STA�u���q��uNC�s1=�� C��o'��|,d�_ m��������Ǐُ� ���!�3�E�W�i�{� ������ß՟|+��� ���[�&�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���2� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� ���*�<�N�`�r� ������������ �&�8�J�\�n����� ������������" 4FXj|��� ����0B Tfx������ ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? ��?�?�?�?�? OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_�?f_�_�_�_�_ �_�_�_
oo.o@oRo dovo�o�o�o�o�o�o �o*<r_`r �������� �&�8�J�\�n����� ����ȏڏ����"� XF�X�j�|������� ğ֟�����0�B� T�f�x���������ү ���,��,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������ �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/��/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO �/�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6olOFolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��Ro@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟ޟ�� 8�&�8�J�\�n����� ����ȯگ����"� 4�F�X�j�|������� Ŀֿ����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������ ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������� �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?��?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ x?f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o L_&L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���2 �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ���*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶���������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x��������� ������,�>�P�b� t��������������� (:L^p� ������  $6HZl~�� �����/ /2/ D/V/�f/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�?��?I�$ENETMODE 1>r%��  _   4@4@�<E7OIH@RROR�_PROG %�#J%�LH�OLFdETABLE  #K�|/�O�O�OJRR�SEV_NUM �2B  ��-A)PdA_AUTO_ENB  PE�+CaD_NO>Q �?#KEA(R  �*��P��P��P��P4P+�P�_�_�_ZT�HIS%SLA+@S[_�ALM 1@#K� �LD�\�@+ �_;oMo_oqo�o�o�_�_R`P  #K�QFB�j@TCP_�VER !#J!��O�o$EXTLO�G_REQ�V�QY,sSIZ5'tSkTKRyoU�)r�TOL  LAD�z�R�A 't_BWD�`�pHV�qDww_DI�q Ar%�STDDLAKB�vS�TEP��@�pO�P_DOtbAFD�R_GRP 1B#INQd 	�or�F@�c��[��w���#/[��7u���� �����c����ɍc�C�!C���B[�A���AA�wtA����΍B�ωB��L]B8�?A�9LArKA�aH΍ɏ?�*�c��N���r�����  A��b]A��7>煖���D@
 �K_&�֑Β�C��b��ׄEݐ�F,D :�D�`�E���)�D  Ew�� b�D+�m�{C�(�C��N���B�ƈ��΍@UUU��UU��ۯ&�~8��� E�@����΍OHcGP{)�K��6�/Jk�΍?�R���:G:�z�9{󨂆�΍;n��Į:��|�LA�ϝL�cy�P�E�EATURE� Cr%�pJA�HandlingTool �� svdeE�nglish D�ictionar�y��
! �4D St�ar}d�  ffs���AA Vis� ?Master���� R597�nal�og I/O(� � 90 HS�gle Shift(��R6417�uto� Softwar�e Update�  4 RR��m�atic Bac7kupe�49����ground E�ditI�  oa�diCameKra[�F_�4�t��nrRndIm����duc��omm�@�calib U�I�� ERm�Co�n��@�onito�r��ct\j3�t�r�Reliab�t���PCVL�Data Acq�u=�:���.sv~k�iagnos���X���cflxk�o�cument;�e�weE���'�Ok�u�al Check Safety%�� g H5��hanced Us�гFr���PC��xt. DIO 5��fi�� def.���end��Err�D�L��������sH-����rV��� �p���41m�FCTN_ Menu��v`����H55��FTPw InF�facv�{  J�JG��}pB�k Exc�нg�� Par�T���Proxy S�v��  j616��igh-Spe���Ski� 6.�fd㰎��mmuwnic��ons�������urm�F�_� �R67\���c�onnect 2���04��IncrΈ�str�z�FC�B��KAREL �Cmd. L��u�a��J�Uc�Runw-Ti��Env#��"
c�P�el u+��s��S/W���  �License�Ӳփ��$�Book(Sy�E�m)��! to�MACROs�,��/O3�{��I�F��H���
 8�1 ��MechS�top��t:�z� 7T "j�Mi�w�9 ����Mix��X�����orch��o}du�witch(����o:҉�. d� -��Optm�� R7*���f{il��Pick�zX�g� OAD�?ulti-T�������v
EP?CM funT�z��90#ow�Reg�iE��  d���PnH�t F* D/��[Y�Num Se=l6  ry��y>�� Adju�����k�w�  pr��tatuR*�N�DI��ٵ�r��R�DM Robot>�scove�*�Rem4 �n� �,���	#Servo�� ��?SNPXs b��(�rt ��w�Libr���p#bo��w�� E{ �  m� W o��t�m�ssag P�v��!z�[s in� VC&,Ӧ��` ����(TP�"/�I�� )��� MI�LIB=fxtp~� P Firm���)�d���n�Accd����e�71TXr��L��� eln �<I0� ����ew\mc�1rquu��imulaC��� �te.f�1u� PYa���Ma��T��t^Ѡ&��ev.��~��USB poo V@�iP�a�� ���,@nexcep�t��# n�� �\`@�����n0VC!�1r���:hk�1<��j4<�{+�4<�SP CSUI�к�6�IXC�&ro�Hx��� 
�We�b Pl���97��QC!�Nl21R��@�ԩ�D��3%F� i��gXGrid!play o�gX� ���L� �iRnIVM�Re  e� -2�000iB/16�5��rAscii����1�� 5 (K�UUpl���3�5�s!��!t� rc��Cyct���]�ori��5%FRL��amY*�HMIo Dev�� (Y!����PC��-@o #�asswo&�2
4�9\��64MB �DRA�!	�l2�bFcRO�kY�7�rc�'visD���5c����ell[�L�H54&�sh*q�"�0C|Ac�^�2@Eu��p�6,JDEutyt�s��V�Ict�� .���{ ��sp 2��yaV�B by 
 ���	 B"X�q it�2���T1>�K%.�10�OL�`Su�pB�Rc�OP�T ��njNS �bS�B�cro��c	#<{%�T mjp��='��a�puest*�SuS�`e�tex{�y ���$LimipYb�Sp����1��0�P���gJ�n�Vi�rt��	#���Mdspn�8��h51>oCVIS� IRp�vC�JDIRCALrv>D�+�IC:;0�x ��phicpD�hо�Abui��l�� F�!P�MM�p�� !fl�owh1f.sk�O�SFILE Ar�" u�co gtp���BMON��IX3 c�җ!m T�N@_PTTB:��i���R805� ��J ����
��⊔j�^��m����"PALT=:�`clud����AIW�- Wai�t/Y�ea�� t�k��TP�bDOE�S NOT RE�STO �60Li=n��mark��GuseJ�z ��c�  Synchr@��z���DSUPPR���PRG IN +AR�A ��Ag���OVC_VALU�E�OBLEM ���V��TMi�TM�W��G���ab�A MOTION��STRUCT l���BRAKE �ABNORMx� ���g�$FMS_�GRV0ISMAT�CH=uu�Z�MAS�T HANG U�P 37m�MUL�TI WIN/L�OCB���SERV�O��AG GAR�*�
�GRID D�ETECT BU�A���!0�����TR�ANSLAY�OF� UTX��F� DB/s�DO �PULSE@EN~CCAMERA����c�`REMARK FOR�� w��L�0\h���EX�PANDED POS>���%'�����SCREEl�A�Y CRUSH ��P!�OTN56a0����fԡ�ND�SYRUNNI���Ɛ�USR��F� TOLp�NCEu ��vK�FSE���Ŧ ���S-14w4 A��ART���
p�FA_� CP�MO-073�v�>��ospowᇡ���@�ڢ�ps�ܛЛQ��syde�m�֛б���sno�sv.�Ь��ۛ�i����gA S���HQ�Z�a_cmC�-�PH�T��!  OMRsPA&;6�&`�PR��[qdp�G(Co��Y�P,�" �1�қ��G���<��g�R556����ic��e�|��G��tg��2�G���aHP} ��tplugN�sSp��O�-inb�SPPG ��~�r�C(SC�P`��LC���J�\sw'�� � �� �w��
�^ ����trsv���1�.pc
���  fx�_�2����%3��B	4.:�BB��5���&6�D#�C7�	��B	8���Btn
�0���=��F�n��sN�Nom}i�p Posi�Q����NN�54!9~�Ї�`(B��ܝ���TXP5
no�mpos\nmt�p "NMTX"� #1�П]�e9t6�OMP�.�����-fxuif�N�-fle��b�F�XUFd�Ё�*"(�'�6	"$  f !"*!�sq&_�е�o$�	 ,]�t#w斠rl�o(uf.�vr.��'
@�in�cus.c�o"��#2+1mpmplete"��M?U4 K?]?�?�?�?�?�?�? �?�?�?O#OPOGOYO��O}O�C�p<��A�2�
  �O�O�O�O�O�O,_#_ 5_b_Y_k_�_�_�_�_ �_�_�_�_(oo1o^o Uogo�o�o�o�o�o�o �o�o$-ZQc�}��������� ���
�ya�C7j@���v�t���r�q�j8�47\wti�v ��/���a��/�q���weW ��=���{47,r768R��asyArm&�f�un?�f�C�R� �S01h��Ь�(X�t E����X'��~�\popupcAt�#Ã,��aN��M�-Shelld�R533R��J�/ (Mu��-[����;'���vrdb�c2
5C�%� �enoio.fC�EnH�ced I/Od�"�3���J�6v�ŗ�p��ܷ���repa��c���?�accu�airR�AP�AirS�6;�0�kz� (\�p���O���S��ca
���4�O� �2��!S�� 2 Gu�c�����49 R63z����(������@��g�aΠib�#A�oSEL�^�/����!C�`�n,a�flowL�3� AF-AS-FMS��mmP�AFSM��x�2~勁����(�غ����S�˴��afgl
2��G˾!��P̴ۢF�̳2V�F�e�AFް��������᳣�O/�e�2�ȡ̱��d�̱2NL�AF2�Ͻ�2�� ���l��RӋ1B�@sŚ�w�x���!w��P��G�_�ɶ3��A�!㹽�AS ��~�5� �����`#������LO��.���˱������C�clrpt�hR�w�ic Cl�[���thϜ778ʪ�7��g��ȀBas��@�w��� �ᛲ���>�S��㒐��tpqe=���s�sub����� n��=�� /�w�set��� �"�q���w�A�Off-�line Svu�lari6�>�85x>���[�85 ( ���tya���sia�d\tp� "SIAD�/���x�,k�plug���Dispense� P� j�=�SPL%G. 9s�(����g-i��Q����e�a�\sldsp�i�"�U8���0� }L% Trk F�� ̀<��>��ꖇ%\���For��tq� �(�]tcyc� "T� ���k�tGgtp�/��!l��la��-#ptkmisc5#�"!�����w� ~��os�able EOAT<�_�G�����(@��
� ��3Q!b��"t���%1��Fou���os1�)t�47<�q�47 (U4��on�)0�_�K1�2+3���7�a�J5��r7�0��ervo Tip Dres�F�08>���0ȁ�H7�r7��A\turnd @b���D0�'�����MHb<+�2	��@_��Lq�3�2]?C5/�S��Ai�n`�� �'gch�t ��VG��r�S�GCH J*!J6�43>�Q��GN �CfQ��cT\svosvch��CH/|���TglgouV/�[gnc]���_�P��R�	dV;�sgdi�a�Ssb cor�ey2XDG�P70�P�Q{<�b(~d7�`O8��rc�cinib���x^btdw�j952Ҵ�ut@unSCS<��R Jp�iH8r({��u����q�Pat݂c�w������ux�h86�9I�7�l��

/F,��v��3�� mtsv "M�TSV�X�j983\R���&P�s��ov��&_p���vruk%_c6�� ����pex_�r��col$Q����v�v�"�r���&�sxcM.Tool��k���=MTOF7p84� J571 R8C14�!7E�ǈ�(���q���	mtofs�0��ߘ�2�⒑��pt�a��lletxo���k�PTLC��9����J9�813���H���T�4�9���`k{;��1�a\pmk920 "K�� �S!R����1�Ȥ<����2¢2�_�ި4@���!�ڣ�a6�1¡4��0����E�ܣ�q8�4f�4C�c&0��5f�����ݤ 9�7bf�7C��ަgr@?"GRIP".������1i "OPT�IC��1ݧpalf? "PALF�Q x@�{ĻPSSUC��F!ަcpt "UNcIT�S7mަxf��XFER��ԃ��et��L�U�&ʾŏ>��psysdj���/����mޤopti���Kޥ����7߹�ssu��+�ޤcpG!W�F��er��S�N�t�����sӸ��d+�[�ad�pՂzaAdapt� CtrlF�3q5	0E�G0汫�_�>��l\apa��.��C����a�1l"�g;ui� GUI��T���c[�c��x�ogJoU et+ra�&��u���386F�� (���1r6��re��3��ETN;����X���5x��j72�2\cust_wcv6�R��v7x߈RS�[8�;QU	9x�KUwv102o>Rwvpat-�<T�ange/;U�h`#C j80�W�eldCondMo���H�JK�#7a�Dq (T���iJ?\atk30e����R�1�{�wm]M3ON�_�0\�$� _��$Xg��p��b��"At��%stop�/rù�Ѐ�Zd��y8N4Ci}r��ld Pr���XvF�ׁ��K��1µ�cS7�O1�1\�q�-\?8�at_u�frm.� #ER�7�xcArc Abnvr�l \itob�9  H�552}�121 �[prc��2 �a�1AAVM� ��20 ���J614��@TUP mch "#@�545�PC#B6���VCAM �awam�0CRI9Me_@UIF��#A�28 0`vr_@N�RE�b.@R631��s�0SCH���DOCV lis=i
@DCSUE�#A�045pR51�EIOCe t��05�42}�R�A96 �pC
@ESET ��c
@J5K@��#@�7K@;bMAS�K acryv@P�RXY cw1wB7�%��0OCO Ph�t�B3�s;B2  tQ�B0�p pa#A�@4�;A39�0Fo�@H^SI�LC�HK�@59�@OP�LG ��;A03 <��PHCR :�P?CSP  GW�R36 ��;A54��P�DSW@_f�0M�D;P "FO�@OqP;P�PPRO!���B7 mforkz�B0�UPCMF	e:�@4f507�U�@�5-hg��!fRSTv-f69`clmP�FRD@�SRMC�N	eH930�eS�NBA�USHLB�	eSM�`mextue�B6�fPVC-gq2�`��~QTCP�U�TMIL	f789�5@ups�`PAC��fPTX	eTELUNrd�R9Ef8@�w1 mpush�#@958Ef957�	eUECKYuUF�R�fVCCM	eVwCOR	�k.vS@gIPLU�@I ��{_f�qXC kZ��_@VVF ��WEBP Y��aT�P��t.�pR62�6 T InpCuG�pnF�I=�u ��6�PGS�R�3_q95 718{ P�0738 f�|�1�@
  ��A�C`6�A63 79�4�B523�5R6�5�1Sua553� ��A4�@gC=@1�qED064 ta�mapF���O�6� sths._@L�IO ��w^p��5� - HefPCM�SC��ӂP��51>@STYL t�_@�TOP ��PR5�{@Wave,�PRgSR ��A801U�OL�Ph� v@OP�ISY0��`� wD.��0L�p}��S���t^pETS�f{un�0SLMTY0|��B9 623�Az�`E�5FVRC�0<_��NL tj�wp'001E��2E��93)E��6 j��:@#U0'@BDݐ5MEݐg8 a֐��U0�` 6������5��J?@s@S���0F�361�=�3 ��;�6�@69�U5`*�2faF�_�7 ��݁Za�8Y�04^�9��H_�_PT�up��20dw0��6u���7 ��L�@��8 �"��9u�+us�0U�1aw��`��{@Ʀ�@Ҧ33ݧ138`���`
�@�?7 R.$M��/��K ���9���4i0E[�1̀Se�@
]�2��Ea��1�4��334������zn�e��Roboz��net�������9��!��j>��\srvo��4��@h���x����S�rv�t ROB*:PM'�e��5��G��n�r�b*��ite��ӿ�5�-�̝6�35v��56�4��7@Main>��tatio����6���������o4���S��, '������\��\cc~�� "TORC�������L��cr�V�CR����5>'�xk965��@���N��MО�6�0���;���o_��w5���0ch��y6���Cv.j�k��iw2 ��
��x5����2.���n���3�V�h�z��5���uSif����c�_�3E@H�,�l�����"T�1���T�2�(�Z�l�4z���?������/�l_i��}3�����0� t{���
  Y2�?�jog\dju�i���og��awWmfr� f��F� �ius�� Eq LibJ��6K񄐞S��/3�� (�bA,��2�7�_5'�\�<�� "MF����d5a��n7y57eM��m K��߽Ҡm���g ����̞A�tw1������tw���#���6 'ink��0LR .ќ�6��J852���J�597�98�88�J�!�1^%N6���b�GN �k\etl�@.�CO���O#|A` "ALNK
�>�%rd_�PB�� �"\wr*1O="�"lS ��P$d�S��88����PN A;RC��PRM�3��@B0��N���!8^�<���1SU P��$P��Ç�H���0��|pм3mpana/'p�ȣ0�1�H57X��85n������ �0K�BH@�<��1��bel������R��<D41�HDY�dhen��8<A���D���Cm���EN������D.��E��<�!� kemp��Dh¼3�m:re��2��pEf"sFMIG6�A00��37JR��|P�!�IGC (�P�.�E�%�чߑT� a;vs��IGE��Gџmigco`'�m�n&NA�ц�fa�vavtj�VTP�o/lfrm "S؆pGoYmsy�ASY�qo/lpdhV�PDyH�oYktpdl7�DL�o/lrf�`CRF�d�y�p8�3b:�s�`.vr3h1y�rLO5ccr��p �4c�§��q�@�����������R�RB�Sg�S����.�o���.��Z=fArbt\��`c.2  �w� ���a�b���! TertiB
ELS�P�2�U�g�YL (Co�mmyle s�eU�%)��bգ�s���'�ps01 "�PS��.#le\pscol���u.�6��ry�Pr: ���vׁ�Q�4syrs�r��-���ice Requ��g%���SRS�2K�9�P6k45.�9R S�"H|����(���vb�Ы/�,M�ۂfO� " ��s�O��sr������aP5A��+�m8���2813�P�49Z�89���A��{��Z�.���g�st�M�\����|�8
?�M�utl�v��'�&Q�N����q s�pdramj�!�peed.�pf%�Q���NN05���J67��2NĻ�� j�(�d� RH�-�	D��b ?"RMTX"��Ə~E�  ;�2 "S�0q�Q�D���slmt�o�ft� mi��SmL��H6Q64봷H62F�20�6c07B��P�38e��2 Hk�e�s�;�5�l�62K�79��7�95�79��60U9j�1F�1x�4��e5��2����H6���843[�2s�8215j��6�MT+�"�@��6����f�� "����S��\Af봆봖�0n��- Positi5o�l��esf �F�1N1h�ݻP(���ti��,봥�ǀ�ņn1Z�POS�s� �0� �h�873�r�riv�e Axes+�H�8��4di��(D�ual Dr�sHΕ�Ȅp��C�\B��j�.�kŔ*�ex�sj� De)�1��63����AM Indexjź��x�&�\ami:�s� �mi&�8�c�a�sC��nt Aongle+�CO;�p���봗#COM��Mom�������Ϋ�gou���! ̂�
fl���Envi� m���6k�d��820)����flx(�2� t��r��ionΓ{�ǅK�r772\ic�P�$	� �x0Z˱t;��2atzn������c�TJ�ync�Ins�p��R76��� �#���Xj�r#mSB����T�b5=mK�masyA`j�ܢ�nc\��MA�SIr�{��b�as��ulti-!A�`�6V��7v!� +��5k�NN�P ���se��!\��FGRLK��v�k��hdzՎF봅"fr�lk��&�m
ŊTr4���C��il/-&�e��r7��0Zo�nd ��:���� "ICRZp�%Q�g8�Piabic.]T�IAB0c���0o�e�I�0V�E �0��1 (�1�4���0濡�0�C�2\i�0t� IA˱�����"�@AiciAC@�0b��!�1�1��!�0omain�sDP�1�n C7`[��0e�DLPV�2�0��hpV��P M_@��̘ ��O]B�ưI:A��Єdp�CD�O�F"�0N>I�A�B���0_�Fd%4�e�o@nn Stan��A[�'"� MCNl�>�90�096:��s�5j��0�Q=���H��0���Q�2~Q(Re�m^PkAeSdard�I0��W2�NQ�0\t�prcmuǰCM�U�0Fv��d��SRP\rc�0�q��jBRSUF�173 �0uipp��[��Ae�J61S �59Q�I�0taV"i Eq[A��Ζ�Rǅd�!ȡjt`�Pcp�����Esr��A�Qvb2� �Qi�ha�@xa �0#�-���1 �a:���1 awmgenyl�q�0ener���Weld zQib�oX�0AWMG�U7{o _q(G>t�A�`%�b�;�d�60t[A3r�t�1.y�R msh�cq@�3��n sh�e�qqGR��1CMSC�U�A���RhjQ�(���p�0l�0rd$�1F�8 p[a��u\q�sh� PSH���� X  ������0
   ;(L r wKq�1K/Fe$�Q7�Ij��w\cl
A "J�����0 H\j�Qcle��"E�S�HeӄuybU��`{A�ybmdprm"�8�zali_varsS�<���iconu���dbg"��0Iz�ց?rgpged"��1l�&��� Ԅm_�0�1�i�Q҃m102<؟�e_no��ȕ�wrspq����wrpirS�[q>��0�gas��Y��1��_�s���wr������fyfӯE�inch30|U���extwd����wrc����'�DՂrdS�Q�D�0!�i�����aN� bo���0�Ə(�/i@��RF�p
q���saj��ca��ntKCMAP ���O D�B�)��T�f�ap"Qj�AP�C��Z���0stmN(PSTM.Q{� ��apcevre*a�o��in
Au7a*a��is
�rbCIS�D G�QMete0/`�3�0T56��i�<�cQ��Q7�ar �>�,KQ�Y��(�\sl(�gr0S�14�e���q�	B..i�A������d��/�[a��>ֻ1���Q�d+Q�G 
�(5ф�M�Q�O K�џ� `+�2�`KQ�����B ��Kq��GT��sU�0���0S30le Ac	t�C�8R��Y
AQ�4.��1�㵏�I��-\J�ds��SU^� %����{A�#���s�!�j691.f�1S�ervoTorc�h9��6Jv�K� 91 (�K�A���Q�svt��VR��AsRC
�es4 F���Q4��MU�dq�v�z�vt/���5�+Q tFEv� ՛0"S`���0h for A�lumi��982Λ� 82������; ���a֞�d�L{���oo�q��l���L�ϊ��\srvt.vK�3e��0�0hP�AS`�� A��<^
�S016F�8a(�0�*�(!ez���hS�ATNQ���h`
�"P�QNG���	��2w�ADW����t��ҋ�М�wenmr�8sn�hanced M;ir�bmag ��b7R69�Q90�+�E.'KQ I>!��I�""\mjQr�MI)R�c;� � e$!.b�06b"%�tmbuswtcpy�Mod� / TCP��REˑX nvkAd�8���!K3CP>� \�$�P}m:1"MBUI2���i2d0� i�+�%���p�930�sPRO_FINET��OJ���J93+� �0 (�5��>鋁Y�3�P?pnio ":���x�1"P�q(@RIO��/ǖ$A��u�3)tj#96Od:��@gT�UHc67J�O��Q�`FSW䑡@���?K�67\fswpr��W+F�}�A\f_��ach޷	�A;be�r4���96�p_f�wd!6���f_r�ea/T[O 'Qneu4��_�Rr��sR��C�Qurn���%S�enא� $Ssw��t�_fswcol�#�n�AQ��Ak��cvvcuZ�2�i�RCalib V~z!nc Utl4�OVCUT� ��1?��b(�a��VisF�u�cj���`k�vc�cU���c�tpfia�_z��`p6b�_8+�apset�3���c\z_�p{���k���uKA4���c��j9�88/�To��orYs1�!�p.�=8�?5 �p ^ol +!p��+��p\gf*��D�sT�c���V�Mas@��9�;� �t�ۮ���1� P�osiZ�����or�dt���v�
�02\���up޶�����r�_dc1$AB�As.��I[\N�bj An�e��b���򾿀��ۿ]���+�ޘ�� �_wQW�� k_Bc0y�t{G���F4�1�k�nifi3 sSpeY��94� a�1�UI n���v�>��k1��`�\frco���
�j9��1�Brake ch:ѡf�`0�{Q�5GJ��(�ck�rpȺ���˕51��b��BRCHUCD ����P�����5/�C����m�ulaneous��=���>55`�lo�H�SiɀS�TD u�LA�NG ��!�c�s��0C�T��\�cscsm���1ﳔsﳠ�=��C8ﳡ�N�dss' �Σ@c S�F�
������3�V68��F�,��sﳥ�s\��u�ߣ�ć��N�r69����gn�ost�eo� n������1�U�i -��9��C�ﳵ�7�z!�\�"DVMV����"r6�Đ�ﴃ! !��p��Uԧ� tr�D!ﳢ��2ﳡ�[�4� TcԦ���er�!��q>+�\pc3j��׸��Ƴ075.�os.Re���rN��� g��2c�6��ė�� �|����75\pt�TJC6���b���Ā���Bg�ė@I�>�S�i>��80��J979a�08� 1���(Iepi{�UL+�oﳔ#��a��f "NRU���¡�prsta�2�£��gutl.��RBT��OPTN�q0\?�r?V�@H nr?�ro�vq?l rb?r�DPN���!�r�rdfi���u𷁟�basi1c�ߡ�fc� ��J��A-�q��H�829V �$��9��@������Ph>�c "F2���29���j83���ce C�t�our� UPDT�3�5����Fo��on���aг�Ӵ�Q8�ho�ff���r� 35�fnV���r��\f�V�����\fcn��rg%3($��% ��r�A������6�%�D �E������g0@=��$���$n���/1!46%u��C/ T0\> ](\��0R2��p�0ޖ�0v�0�2v 6`�0���0?U8�0�1�Br�0���0�4U0L�vpofs`1|��1�3>y0� mgp�s�?��6un�Q�,x/@�4s�e�5ҌBT0��b �cellf�1��e�l/@Cp���1��Rp�1�f�B��519�1ll F�B/@��p�/@b�C�Bn/@fncl��"RA��Z/@<^V�Bfndru��AsIND"�1�>�A.�1\fn��t�A^f`/@t�B&PTPexjA �?�@/@%QTPc�1�vp�1u�B&Ptqd~_��[ Q�2�V�Gj7��/@- V-50�0i//@10i 3D�/@�[S��1�5�`ab`�13D�E�/@N��<9\ca�lc@�_.27/@vsfit3Ep/@�{a��/@7�u/@`�`�Tra/@B��KJ�a�MJ�`�b�e�1�b@E��1�/@Ov/@j�`\que�1�?�3Ar�po��8_�`8�1eopush3�� ��$/@}s\�М�v��/��qkm�1ޕ\�swqa�?�h�qainj|wkclb*O��?q�vs
AJ\udsbclt���eenn��g�|wigchk4��uv�avuA�s��� t��6�
  �тv��3��_p��FA��GAv"73�1cro��4��,�v�Apo �/@��8�a�jB��iR��qon Erro�9���.m�FQ�A7�57�Aж�1�� (#iR�A���R.]kZ��<d\mherh�d�AH4P���}��\�ire:AR���r�ee���/0�B@���l4��Z�h:Ahd��� `������j��cv�a����`�1SP AP�AS�A��SASz�0�9 �q CTAM\ڠQTABڡP�AGz�13�Ҷ�Π(�`�Q����p&u/Mޤ�pas\�aama�s+�=�
AF��c��s��bia�B?�����VS����VSI�AС��D�q����(��A��vA8D��  �6� ���
��1  !�   ��� ���/@(�8 ���\���ұ(H��s ��]ia\ia�`�a�`���P��g�QoiZĳ|c�x�����  �����*SYST��EM/@A �����$ˢ�S � �/@��������AT�STKSIZ������/@������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy�� �����	- ?Qcu���� ���*�Ȳ���TART_T �SAG��$D��I�GNAL��SAR�TUP_CNfQ /a/s/�/�/�/�/�/��DK�2!
�
 �/??)?;?M?�_?q?�?�?�?�?�:�99�@L���$FEAT_DE�MO C�����1@   �8MO OMODO VO�OzO�O�O�O�O�O �O_
__I_@_R__ v_�_�_�_�_�_�_o ooEo<oNo{oro�o �o�o�o�o�o A8Jwn��� ������=�4� F�s�j�|�������̏ ֏����9�0�B�o� f�x�������ȟҟ�� ���5�,�>�k�b�t� ������įί���� 1�(�:�g�^�p����� ����ʿ��� �-�$� 6�c�Z�lϙϐϢϼ� ��������)� �2�_� V�hߕߌߞ߸����� ����%��.�[�R�d� ������������ !��*�W�N�`����� ������������ &SJ\���� ����"O FX�|���� ��///K/B/T/ �/x/�/�/�/�/�/�/ ???G?>?P?}?t? �?�?�?�?�?�?OO OCO:OLOyOpO�O�O �O�O�O�O	_ __?_ 6_H_u_l_~_�_�_�_ �_�_o�_o;o2oDo qohozo�o�o�o�o�o �o
7.@md v������� �3�*�<�i�`�r��� ��Ï��̏�����/� &�8�e�\�n������� ��ȟ�����+�"�4� a�X�j���������į ����'��0�]�T� f������������� ��#��,�Y�P�b�|� �ϳϪϼ�������� �(�U�L�^�x߂߯� �߸���������$� Q�H�Z�t�~���� �������� �M�D� V�p�z����������� ��
I@Rl v������ E<Nhr� �����/// A/8/J/d/n/�/�/�/ �/�/�/?�/?=?4? F?`?j?�?�?�?�?�? �?O�?O9O0OBO\O fO�O�O�O�O�O�O�O �O_5_,_>_X_b_�_ �_�_�_�_�_�_�_o 1o(o:oTo^o�o�o�o �o�o�o�o�o -$ 6PZ�~��� ����)� �2�L� V���z�������� ���%��.�H�R�� v������������� !��*�D�N�{�r��� �������ޯ��� &�@�J�w�n������� ���ڿ���"�<� F�s�j�|ϩϠϲ��� �������8�B�o� f�xߥߜ߮������� ���4�>�k�b�t� ������������ �0�:�g�^�p����� ��������	 , 6cZl���� ���(2_ Vh������ /�
/$/./[/R/d/ �/�/�/�/�/�/�/�/ ? ?*?W?N?`?�?�? �?�?�?�?�?�?OO &OSOJO\O�O�O�O�O �O�O�O�O�O_"_O_ F_X_�_|_�_�_�_�_ �_�_�_ooKoBoTo �oxo�o�o�o�o�o�o �oG>P}t �������� �C�:�L�y�p����� �����܏���?� 6�H�u�l�~������� �؟���;�2�D� q�h�z�������ݯԯ � �
�7�.�@�m�d��v�������ٿп��  ��$�6� H�Z�l�~ϐϢϴ��� ������� �2�D�V� h�zߌߞ߰������� ��
��.�@�R�d�v� ������������ �*�<�N�`�r����� ����������& 8J\n���� ����"4F Xj|����� ��//0/B/T/f/ x/�/�/�/�/�/�/�/ ??,?>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^OpO�O�O�O �O�O�O�O __$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�o�o�o�o �o
.@Rdv �������� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�F� X�j�|�������į֯ �����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ������� *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�?|�?�9  �8 �1O(O:OLO^OpO�O �O�O�O�O�O�O __ $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p��� ������������  $6HZl~�� ����� 2 DVhz���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�?�?A@�8O,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o  2DVhz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�xϊϜϮ��� ��������,�>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� � �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿����$FEAT_�DEMOIN  �Ā2������INDEX'��6���ILECO�MP D���h�5��^��SETUP2 �Eh�r�� � N ��[�_AP2BCK 1Fh�?  �)���"��%�����k��� /����[����ߌ� ��D���h�����3� ��W�i��ߍ����� R���v�����A��� e������*���N��� ������=O��s �&��\�� '�K�o� �4��j��#/ �0/Y/�}//�/�/ B/�/f/�/?�/1?�/ U?g?�/�??�?>?�? �?t?	O�?-O?O�?cO �?�O�O(O�OLO�O�O �O_�O;_�OH_q_ _ �_$_�_�_Z_�_~_o %o�_Io�_mooo�o�2o�oVo�o�owɫ�P�� 2��*.cVRN�`*Q�w�c}��e8pPC����`FR6:D��~�"��{TF� F�X��uC���)�����f*.F;ُ�a	�sǏ���*���STM J�S�^��p�K����`iPe�ndant Pa'nel����H����p�ϟ���3���GIF=�g�r�S��"�����JPG���r�ׯ0����;��zJSE�n��`�\��%
J�avaScript��ůCS���q��߿�� %Cas�cading S�tyle She�etsϐ`
AR�GNAME.DTMϰlu�\a�ρ���Ģ�N�	PANE3L1����%u���%ߜ�����2߀�� n�+�=�����3���@��߯���V���4"��v�3�E���Y�T�PEINS.XML��}�:\������Custom T?oolbar6��h�PASSWOR�D��nFRS:�\y�8� %Pa�ssword Config���o ����9�o]���� "�F��|� 5��k��� �T�x//�C/ �g/y//�/,/�/P/ b/�/�/?�/?Q?�/ u??�?�?:?�?^?�? O�?)O�?MO�?�?�O O�O6O�O�OlO_�O %_7_�O[_�O_�_ _ �_D_�_h_z_o�_3o �_,oio�_�oo�o�o Ro�ovo�oA�o e�o�*�N� ����=�O��s� �����8�͏\�񏀏 ��'���K�ڏD���� ��4�ɟ۟j�����#� 5�ğY��}����� B�ׯf�Я���1��� U�g����������P� �t�	Ϙ���?�οc� �\ϙ�(Ͻ�L����� ��ߦ�;�M���q� � ��$�6���Z���~��� %��I���m���� 2�����h����!��� ��W���{�
�t���@� ��d�����/��S e����<N����$FILE_�DGBCK 1F���� ��� ( �)�
SUMMARY�.DG��MD�:!a� Di�ag Summa�rybo

CONSLOGW:L���tConso?le log�n	TPACCN��@/%(/e/pTP� Account�in/o
FR6�:IPKDMP.'ZIP�/�
�/�/�q� Except�ion�/�+MME?MCHECK[/��Pq?�Memory Datar?�ra,])]1HADOWg?L?^?�?��3Shadow� Changes��?�-��)	FTP�MO�?QO|7��mment �TBDzOr=t�)ETHERNEToO�01�O�Ot�Etherne�t �figur�a?udADCSV�RFnOTOfO_�1�%DP veri?fy all�_��10"�?UDIF�Fw_]_o_o�0%=�Xdiffo�W|01DPCHGD1�_8�_�_�o o�o�S!�Gi2ofoxo� �o4�oG�D3�o�o� �#�GvUPDATES.�p��?FRS:\���uUpdate?s List���PSRBWLD.CME���Y����PS_ROBOWEL�Omޏ��� ��8�J�ُn����� !���ȟW��{���"� ��F�՟j�|����/� į֯e��������� T��x������=�ҿ a���ϗ�,ϻ�P�b� ��Ϫ�9ϣ���o� ߓ��:���^��ς� ��#߸�G�����}�� ��6���/�l��ߐ�� ����U���y�� ��� D���h�z�	���-��� Q���������-R ��v��;�_ ��*�N�G ��7��m/ �&/8/�\/��/�/ !/�/E/�/i/�/?�/ 4?�/E?j?�/�??�? �?S?�?w?OO�?BO �?fO�?_O�O+O�OOO �O�O�O_�O>_P_�O�t__�_�_  �$�FILE_�PR�����P�����XMDONLY 1F�U~�P 
 �;_ o__6o�_Colo5_�o o�o�oUo�oyo  �oD�ohz	�- �Q�����@� R��v������;�Џ _�����*���N�ݏ [������7�̟ޟm� ���&�8�ǟ\�럀� ��!���E�گi���~�ZVISBCK�X|�Q�S*.VD�|a�ϠFR:\0��ION\DATA�\L��ϠVi�sion VD file����տ� �����/Ͼ�@�e��� ��ϭϿ�N���r�� �Ϩ�=���a�s�.ߗ� &߻�J����߀��� 9�K���o��ߓ�"�4� ��X������#���G� ��X�}����0����� f���������U�Z�MR2_GRP �1G�[�C4�  B�> 	 ��Q��� E�� E�@���`
� OHcGP��K���Jkǅ�?� `� :�G:�<9{��<H�A�  dv{BH�C��N�OB�ƈ�`�}� z  D����>��	@UUU��UU�`/����#@=udѽ���H=��=�~�=�yC,����;�.;�!�9���:�b:�l?���/ /�/�/�E� � F,D �!D��`�#�u�-��E��� �!D+�2C��dR_CFG {H�[T �/�O?a?s?�NO ��X�
F0��1 �0 �  ���0��PRM_CHKTYP  �P��> �P�P�P��1O=M�0_MIN�0<g���0�PX�P�SSB%3I�U�P�#O:CCO�UO�UTP_DEF'_OW�P:�YpA�IRCOM�0{O��$GENOVRD�_DO�6�R�LT[HR�6 d�Ed�Do_ENB�O �@/RAVCxJGC� ��[OF_�/j_��x_�_7�P��QOU{ P��B�8��(�_�_�_oo  C�f`\Vo�X�oYm%~oBȽ�b�	�Y\\OPSMTSQY�� @ed�$HOS�TC%21R9�[�G 	;x;{�;8k�ye������z���1�C�U�xy��	�anonymous|�����Ώ��7: L^3�r���{��� ���� �՟����� @�~���e�w������� ��� ���4��h�=� O�a�s�������Ϳ ߿��R�'�9�K�]� oϾ�Я⯈�����*� ���#�5�G���k�}� �ߡ����������� �1�ϒϤ϶ϸߝ� ����������	�X�-� ?�Q�c���t��߫��� ������B�T�f�x�z� _������� �%7Z��m ���(: <!/pE/W/i/{/�/ ��/�/�/�/�//Z lA?S?e?w?��� ��/�?2/OO+O=O OO�/sO�O�O�O�O�? ?.?__'_9_�mq�ENT 1S�[� P!�O�_�R  w_�_�_�_�_�_�_ o �_,ooUozo=o�oao �o�o�o�o
�o�o@ d'�K�o� ����*��N�� G���s���k�̏���� ����׏%�J��n�1� ��U���y�ڟ������ӟ4���X��QUICC0e�A�S����w�1�������w�2����T�!ROUTERU�1�C���!PCJOG�����!192.�168.0.10�~�s�CAMPRT,��ѿ!�1���RTn� �2ϓ�YTNAME !fZ?!ROBOϛ��S_CFG 1R�fY ��Auto-sta�rted�4FTP�?,��?�OW��? {ߍߟ߱���hO���� ��@�.���e�w�� ���6��)���=� _��F�X�j�|�K�� �����������0 BTfx�?�?�?� ���3�,> bt����O� �//(/:/��� �/��/��/�/�/ ? ��/6?H?Z?l?�/�? #?�?�?�?�?�?K/]/ o/O�?hO�/�O�O�O �O�O�?�O
__._QO R_�Ov_�_�_�_�_O O1OCOE_*oyONo`o ro�o�oe_�o�o�o�o o�o�o8J\n� �_�_�_o�;o� "�4�F�X�'|����� ��ď�i�����0� B�����ɏ��� ҟ������>�P� b�t�����+���ί������T_ERR� T���"�PDUSIZ  ���^ɐ�9�>R�W�RD ?�Ō���  guest��������ȿ�ڿ쿣�SCD_GROUP 2U�̫ ����1��!x��2�ǒ  ,C��	$SVMTR_�ID 2�Ti��$GRP_2�$�AXIS_NUM� Y�z�f�NF���SV_PARA�Miɑ� ,$�MOT_S��TT�P_AUTH 1�V1� <!i?Pendan����Jũ���!KAREL:*��݇KC3�C�U�+��VISION SCET��ߊ���!�� ����(������e��<�N��r����CT_RL W1������
��FFF�9E3�FR�S:DEFAUL�T�FANU�C Web Se/rver�
��z� ���������������� �WR_CONF�IG X!��m��"�IDL_CPU_PC0����BȊ�K  BH1MIN<)�OGNh�O+�`���7��3 NP��IM_D�O��TPMO_DNTOL� �_PRTY�K�OLNK 1Y1���#5GYk|}�MASTE� ����	OSLAV�E Z1����O�_CFG��UO�����CYCLE���*�_ASG s1[l�
  ]/o/�/�/�/�/�/�/ �/�/?#?5?G?�0"ď�`�5�_��IP�CH/���RTR�Y_CN0���SCRN_UPD_���9� ����\1�&�O&��$J�23_DSP_E�NB�01�%�@OB�PROC%C��J�OG�1]1��8��d8�?�R;�OR??U�S��LQ�O�O_#_�OG_Y_�k_}_��'ҟ_[CP�OSREEO�KA/NJI_�K��S$1��3^���U�_�UCL_L[ m2�?��PEYLOGGI�N�&��}A9���$LANGUA�GE m��2*� �a"�LG�2�¬������x&аҘP���Q ���'0ꩨ����MC�:\RSCH\0�0\�}`N_DISP `1�����8�O�O �LOC�B�Dzj�A�cOGBOOK a;+�~@����q�q�pXCy�����*�b=�0�O���	�u��y��Fu����!ua@B�UFF 1b ��2��ڏ�r���� ���$�Q�H�Z���~� ������Ɵ������ �M�D�V�����DC�S d�} =���L�����!������!���IO 1e�;+ 
OZ���� Z�j�|�������Ŀֿ �����2�B�T�f� zϊϜϮ����������
�5�Ez TM  2{d�_c�u߇ߙ� �߽���������)� ;�M�_�q�����8��qw8�SEV�02}]4�TYP@�R�`3�E�W���QRS? �Ko���2FL 1fC��0�˯������`%7h�TP_`�@�"�k}NGN�AM%D�e���UP�S*pGI�5a�5��_LOADB@G� %2z%MA�NUTENTIO�ND�MAXUALRMm7�{8�'_PR�4�0�sM�C-pg;)[�q�s�Pc@P 2h�V ��	"���0���t�� ��� /ɨ/O/:/ s/V/h/�/�/�/�/�/ ?�/'??K?.?@?�? l?�?�?�?�?�?�?�? #OOOYODO}OhO�O �O�O�O�O�O�O�O1_ _U_@_y_�_n_�_�_ �_�_�_	o�_-ooQo coFo�oro�o�o�o�o �o�o);_J �fx��������7�"�[�D_LDXDISA� �B�3�MEMO_A�P� E ?��
 �c���ɏۏ�����#�5�IS�C 1i�� � M����b����L�՟�����J�C_MST�R j���SC/D 1k����g� 韋�v�����ӯ��Я 	���-��Q�<�u�`� ������Ͽ���޿� �;�&�8�q�\ϕπ� �Ϥ����������7� "�[�F��jߣߎߠ� ��������!��E�0� U�{�f�������� ������A�,�e�P� ��t��������������+O:s	�MKCFG l'��n�LTARM_*�m���q���,METP�U9d��/�ND�CMNTd�% � n'�c���{�%POSC�F1<PRPM�0�STOL 1�o'� 4@C�<#�
�n�/' �//1/s/U/g/�/ �/�/�/�/�/?�/	?�K?-???�?k1%SI�NG_CHK  y�t�ODAQ��p�=���5DEV� 	'�	MC}:�<HSIZE���C�Ȼ5TASK �%'�%$123456789 \O�nE�7TRIG 1	q`��%H��OA��O0�O�O)�>FYP)A�E��4�3EM_IN�F 1r�� `)AT?&FV0E0�Og]�)OQE0V1&�A3&B1&D2�&S0&C1S0}=V])ATZg_�_�TH�_�_vQ�Oo�XAo?o�_coJo�o�o M_�oq_�_�_�_ �_<so`r%o� Q�����o�o&� �o�o�on�y3��� ȏ�������"�	�F� X��|�/�A�S�e�֟ ����1��0��T�� x���q���a�s�䯗� ����,�>��b����� A�K���w��ǿ�� ɯ:�����#���G� ������ϡ����#��H�/�l��?NITO�RLG ?K  � 	EXEC�1j��2��3��4���5��@��7��8
��9j��6��� ������������ �����������2!�2-�29�2�E�2Q�2]�2i�2�u�2��2��3!�3�-�3�һ1R_GRP_SV 1s<[� (s1���G��I�ܽXͧ�k��Im���n�=FA_D�,N��PL_NAME �!S���!�Default �Personal�ity (fro�m FD) �R�R23� 1t)4?�x)4�����0@ dp* <N`r���� ���&8J\n�82����� ���
//./@/�2<�j/|/�/�/�/�/��/�/�/??0?B? �  �\  �  ��`���  A�  BUm0Tm0��0
Y0��]0����  �Y�i0h0Bm0pm0o�  C�0C�0�P D�  D;���2E@�2�2z�0�1�0�1�2�0�9��2�0�6�4EK  E+� E��6��2�0�2 A DJZ� �3A@DI�2�5�4�9�:�1;�7�:�5�@�5@�O�;�O�3�1�1E�1���0�` E��\�G�4E���C�@ Q�A] Y$UP�5#V��DQL]hT�FQ8@ �B UA U�T�R YU Q|UU�@�Y�Q�] �Q�Y�@B�YAP�1 �R4oBg�UXo�S�1Q `ong�Q�o�o�o�W�o �o�o 2DV`t�U0E	��E�á�orT1T1O�  !l0��{q�d�s�t ��y���tpI<Z*d����y����`q�0 b�[T� @�5?h0�p�T�?q�p�q�@uþ�5o���;��	l��	  ����p�XJ�����X � � ��, �ނO�K���K�zK��ɜK@0>KH?�K$�����О����5��N�?�{�P�@'�6\�����"��Iڿ��
��}v�����X�������0�
�=ô�0�0��� � >ڃ���#�^���l�Y"�0 ��q����͔��'���h������  �T��  ��`��v��	'�� � ��I�� �  ��-`�:�È��ß�=���إ$�@���Z����BZ��t'�5�o�N��j�  '��O�@���?��@�t�@��@����X���MBd0Cf�0��B�1���q��C%���V�/ � W ��^�/�AB-`���$Ń��� ��A�q��1ș_φ�o�p�πϹ� �
�`�����n� �x��ݱ�� ؀��:�m�����?�f�f��0��� ���d�v�%��ߛ�?KY����|��(q���P�����ȃȄ2��?33�������;���;���;��D�;�$;�< Jl ��=�L�~�Z���=�?offf?��?&z�ޡ�A���@�,��j��u၄�� p���n���^約O�$� �H�3�l�W���{���`������+���F�p ��&��J��k��=,�ɘD�@����0�  F���� ��5 YDV �z�ƚG���/ a'/�N/�r/�/�/4�/G�A�0����O�tp��B�0h/?d/%? ?I?4?���pA�0t2 -`|1�?�u�?\?�2;�<��Ŝ?���?�?hOO*�į��W*O�C��@�` Ca'O*�4��0�1�A���ܨ���C>�CR BA��Aˉ7࢙���"���z���q��=��\)xO� ʊ=��=qA�B)�{���O� ��(��g�/P�q�Bp���{���8R��K����J?&DK���	HwW�H�'���!��LA�L��9K��4HŀHH� h_�zP��Lm��J�sdHK� ?H-�A��_wO �_�_o�_%ooIo4o moXojo�o�o�o�o�o �o�oE0iT �x������ �/��S�>�w�b��� ����я�������� =�(�:�s�^������� ��ߟʟ�� �9�$� ]�H���l�������ۯ8Ư���G�$��� C���4�F@��8��u�8�V����������Ͽп�����?��F( Q�`���G� ���x�8E��Y��>x�	3Z�q_�Ϧϴª�����ϰ�fC3�g����̅��?�3�Ȭ�ـX�F�|�jߠߎ��5P��P������N�`����.���P�0b����7���
C@�C@5����
� @�.�d�������������������������&  ?JK  �@^���v�����2 wD�J�E����0��B}1q1}0C)�f@�AC@@�?CB�J�J�m��C�����R���3��E�(��F���
/�/**@9$���4�C@C@���4�;
 */�/�/�/�/�/ �/�/??/?A?S?e?�w?�J�2��������$MSKCFMAP  D� �g!c!�>�3ONREwL  s��1��а2EXCFEN�B�7
�3�5AFN�CODJOGOV�LIM�7d@Bd��2KEY�7eE��2RUNULeE��2SFSPDTY���FE�3SIGN|�?DT1MOTWO�A�2_CE_G�RP 1zD�3\,�;_$�__q_� [_�_S_�_w_�_�_�_ o�_oPooto�o=o �oao�o�o�o�o�o :�o^pW�K�������1QZ_�EDIT�D�7�3T�COM_CFG 1{�=r&I�[�m�}
)�_ARC_B���DIUAP_C�PL��(DNOCH�ECK ?�; �������
� �.�@�R�d�v����������П����;NO_WAIT_L�Gl�	PNT1�|�;zi+F�_ERRQs2}�9�ф �����ï���3���^ńT_MOt�~{�x OZ��D��8�?�_�I��b 6�m�PARAM:u��;�f&4����w� =� 3�45678901 '�9�K�"�j�|�Xψπ���Ϡ��������w��,�>�ѿb�ƃUM_RSPACE�?�R�o��ߥ��$OD�RDSP���F$HO�FFSET_CAqR�����DIS�����PEN_FIL�E��Ao����PT?ION_IOvO�A�;�M_PRG %��%$*t���WORK �W'C ���6���2���S���	� �a���6�C����RG_DSBL'  DCj,@����RIENTTO��0���2 ��UT_SIM_DC���2�2��V��LCT �P�����>��_PEXE���GRAT��\F$E��>��UP ���x E �/A'es	��$��2St)4��x)4����@ dRߺ�� �&8J\n ��������/"/a�2�R/d/v/ �/�/�/�/�/�/�/��<A/?0?B?T?f?x? �?�?�?�?�?�?�?������)P�  ��  �p�A� g B!@�B�Y�@H@�  ���@p�B!@p�!@�d�c���P �D�  D��NbBE@jB_Bzd� `A`@{A{Bx@�I{Bd@��F|DEK  E+� E��F�Bx@0kB�A�D�JZ�fC�A �D�I�B�ElD�I�JlA;eGJ�E<P�Ec_}KPs_aC[A{AEhA�m@?�` E���WxDE���S��@�Q�Q@�]�Y�U�P�E�V��T �Q md�V�Q�@�R�U �A�U@dcb�Y�U�Q0e�U˵@�ida�mda\i <P�B�i�A�P[A�b�o �g�e�chA�Q"w da4Bp�gx�� ����
����"�A @E�W���P�s� ��j�����(�(��� �O 1y(�Ho(�&��`�o0��C @�Eo�o��?|��C@�E��.�  ;��	lo�	�� ����p�X̰��q���X � � ��, �����H����H��H�P�uHV�2H�H_3��<���&��B�!@	�C����@�γ�4@L@�/
=�g��`@D��(�:�L�)�Aß�w½��ªV y�H@����p�ˣQ��֡�hD��D��  �  �������Q�6�%�	�'� � T��I� �  y��`R�=���x���(�@�������ʿ;��$�߯�r'�Np�"�  'F��:ą�Ca�B@CfBd�B�Au�G�Y� ��  ��C%�  ���^
��/V�B�`��p���;� ������wA ���^�'�M�8�qߨ��
�`��U�n� �x������ L����:O���Q��?�ffǏ���� z߶�%�ㅡ8��E�.S�?Y����4�|�	(����P���ő�������?333Q�����;��;����;�D�;��$;�< J!l�����6�޳8����?fff?��?y&2�A�D�@�,P�Q���-� 9�T�(���&����l� ����� ��$H 3l~i���� ��s������V���Dڹ@�U�@�  Fg�D��� ���/�/G/2/ k/�����-]/�/�/ =?y/*?<?N?`?��AL@��j��	�d�B8@ ?�??�?�?O�?B�'�A�*D�`4A ;O�0�?bO����S�}�?�؏O�O�O�O�Q��g��W�OC�>�P�` Ca�O�*�D��@�ALQ@I�	�b���C>�CR BA��Aˉ7��Q���"���z���q��=��\)0_�0ʊ=��=qA��B)�{�녨_�0��(��g��P�q�Bp���{���8R�MK����J?&DK���	HwW�H�'���1�MLA�L��9K��4HŀHH�  o�2`��Lm��J�sdHK� ?H-�A�Jo/_ �o�o�o�o�o�o�o %"[Fj� ������!�� E�0�i�T���x���Ï ���ҏ���/��?� e�P���t�����џ�� �����+��O�:�s� ^�������ͯ���ܯ � �9�$�]�H�Z���8~����KG�$��ſ� C�����@��8?�-��V��7�>�w�b���ψ�r������ϲV(xA�`����ϸ���0��ų�Y«N0߲S3Z�q_L�^�lҪ�x���߰�fC3�g��߶܅��?�3�Ȭ���ـ���4�"�X�F�EP��P��!�/���`�������`���0�S�>�V�7`�r�
{�{5��V����� ��������/I ��JXj�t��̪�����  ?JK  ���@.dR�r�2 wD��E���0�VB5A)A5@C)�P��A��@9O�X/"/2,C����2/�[/i*�CN�E�(�VF�i/�/�/�/R�*@�$�XxD�����O�|D�K
 �/E?W?i?{?�?�? �?�?�?�?�?OO/O�ZB��\������$PARAM�_MENU ?��� � DEFP�ULSE;K	W�AITTMOUTޓKRCV�O �SHELL_W�RK.$CUR_oSTYL�@�L�OPT��OPTB��O�BC�OR_DECSN�@{�N\H_Z_ l_�_�_�_�_�_�_�_��_%o o2oDomohAS�SREL_ID � +�x�@}dUSE�_PROG %�wJ%io�o}cCCR�@+�C�g_HO�ST !wJ!�d#�jT���o?s�qAs{�k_TI�ME�B�f�eh@GDEBUG�`wK}c�GINP_FLM1S�~�xTR��wWPGA � �|N���CH��xTYPEtL� hobo�� ����Ώ��	���(� Q�L�^�p��������� �ܟ� �)�$�6�H� q�l�~�������Ưد����� �I��uWO�RD ?	&�	�RS��PNeS��D��JOQ��TEbpF�TR�ACECTL 1���A ���M e���� ߾��DT Q����ӰD �{ z�
��#�0)�0�-�;�M�_�qσ� �ϧ�9����ϯ���� %��)�[�M��qߣ� ���߹�������!�3� E�W�{�������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G)�_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�S/����ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ��������� +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O��O�O�O_Y�$P�GTRACELE�N  Q  ���P��'V_UP �����VQ^PBQ�WP'Q_CFG �VU@SQgQ���T9P�_�\kRD�EFSPD ��v\Q9P�'PI�NnPTRL ��v]P8�U�QPE�_CONFIrP�>VU�VQ�T��Y'PLIDoS��v]�QEaGRP 1��gP�Q�C%  �ᙚ�QA�=qGY�� GcX Fg@� A�  D	��T	�Pd�T�i�i�5a5`� 	 p�_�R�[�o ´s�o�kBp>q�T>x�rH9B�!����~� �<T��<]/ ����U�@�y�d� �������я��⏠`z�%�P
�M��� ]���n�����˟��� ڟ����I�4�m�X������!Q
V7�.10beta1��V @�p��@z=q@��R|�aʡC  C5P{B|ܣDf@ ��C�`� D��� D� C��`�`B�䠃`C/�`p�R�r�`1��C�U�$�BdKNOW_M  �U~VBd�SV �mi�-e:�ſ׿� z����
�CσR�mAc�Mfc���8Plڢ	<�Rܡ  �b�� ^����S��ˠ`����I�iRLMRfc�Jy�T�z��QCz�`���u8�J�6mSTfa�1 1�V[
 0a-e��$բ�  �� �߽߫�������4�� )�;�M��q����� ���������T�h��2s���Q�<��a�3r�������l�A4��������l�5"4Fl�6_q��l�7����l��8�!3l�MA�D3V ^Vh�PARNUM  V[q2πj�SCH� ^U
�� )@S%UPD���e\/�_CMP_o�3PWP�P'WjS_ER/_CHK�%|X�&�/�+RS�}�Ba_#MO��/�%_�/\e�_RES_GrВv� ��nr?e?�?�? �?�?�?�?�?OO8O�+O\OOO�_44q�>< N?�O35��O�O�O53  �O�O _53^ _:_ ?_53� Z_y_~_53�  �_�_�_53K�_�_�_52V 1�v�$1���@c���"THR_INR0"!W�z(5dkfMASSxo� Z�gMNwo�cM�ON_QUEUE� �v�	6#0/�*�TNy U�!N�f�+��`END�a?yEcXE(u> BE'p|	�cOPTIOw�&;�`PROGRAoM %�j%�`�6o��bTASK_�I�o~OCFG ���o���DA�TArÖ�@0�2��t��������� g������(�ӏL��^�p���5�INFO
r×Q���d=�ڟ� ���"�4�F�X�j�|� ������į֯������0�B������Q� �lI�� DIT �����5�WER�FLIx^ci�RGA�DJ ���AЋ  ��?#0�d�R�G�a��y���?���a�<@���ɖ%ah�ϸ���[2����`\hF�]b2�2�A(dɻt$��*��/�� **:��#0��d��v���������W�Ab5�Ac	� �-�?߬�c�u߇ߙ� �߽�����N�I��)� ;��_�q������ ��������%�7�I� [�m������������ ����!�EWi {�����/� ��Sew� ������// +/U/O/a/s/�/�/�/ �/�/�/�/??'?9?K?]?�? 	 ��?�? O�7��9O��OfOO��O����PREF S�%�OpOp
۵?IORITY�g�}�߱MPDSP�q�Ϳ�GU�g��ڶOG��_TGʰ�r�j*R�TOE�`1���� (!AFs`E��`s_~W!tc�p~_�]!ud��_�^!icmX�_8o+QXYà��;�Oq)� ��2oDoOp�,omoPe\o �o�o�o�o�o�o�o �o;M4qX��	*)Sâ�MU���^��?(!��6��!/���K�V��~ȁ����AG�,  ��@w�������͏�E��t�C��O�Cղ߱PORT_NUMS�����߱_C?ARTREP�@�����SKSTAW �J�SAVE ���	2600/H738҈O�OTr�`������L���7����7Z�URGE_ENBʹ��aWF(�DOV{�EV�WlPI�ձ)�WRU�P_DELAY ����=�R_HOT %�ֲ=�ɯ�Z�R_NORMA�L��򲸯�ܧSE�MI��Q���QS�KIPȓ��� x}O��yO��̿޿�� �=ϱ���4�F�X�� |�jψϲ����Ϝ��� ���0�B��R�T�f� �߮��߆�������� ,�>��b�P���� p�������(�2��$RBTIF7_>�ARCVTM[BT��E�DCRm���t� Э�E�� ��AEQٿ�C��|A����9 �E��� �������A�o��È݅��"3����� ;���;���;��D�;�$;�< Jl��Se ���� �����	-�?Q�GRDIO_TYPE  ϝ�G]EFPOS1� 1���
 x ?��Z@�</�^� �/v/a/�/5/�/Y/ �/}/�/?�/<?�/`? �/�??1?C?}?�?�? O�?&O�?JO�?GO�O O�O?O�OcO�O�O�O �O�OF_1_j__�_)_ �_M_�_�_�_o�_0o��_To��2 1����oJo�oFo�o<jo�3 1��o�o��o�o`K�S4 1�+=w�����S5 1� ������u���,�S6 1�C�U�g�ࡏ�
�C���S7 1�؏���6�����|؟V�S8 1�m�����˟I�4�m��SMASK 1�z� �������XNO�w������MO�TEL�۫��_CFG ��b�����PL_RANG��O�Q�OWER �����#�SM�_DRYPRG �%�%�����T?ART �|�ʺUME_PRO�����&��_EXEC�_ENB  ��W�GSPD��A�IȜ��X�TDBd�v�R�M��v�MT_��T�w��E�OBOT�_ISOLCخ�F�2�b���NAM/E ��É�OB_ORD_N_UM ?|���H738 �~  ����r����y� ��2�Dr�h�z�}�r� ����r�����
r��x�+��PC_TIM�Eg�S�xE�S23�20�1�����L�TEACH PENDANi�,����7���PM�aintenance Cons���$�"��TKOCL/Cٰp�����o� No Use��N��9ߎ��NPO��^����Y���CH_�L�����	�=��MAVAIL�SѸ�K�����SPACE1 2�� �K�����2�ļ�K�L�b���8�?����� IjAz������ ���':�_ pW������ �S'/:/�_ p/W/�/�����/ /#/?6?�/K?l?S? �?�/�/�/�/�/�?? 1?3?�?GOhO?OQO�? �?�?�?�?�OO-O_ }OC_d_v_]_�O�O�O �O�O�__)_o<o�_ a_roYo�o�_�_�_�_ �oo%o8�oMn U��o�o�o�o�o�o �z�I�j�A�� ��������/� !��E�f�x�O�a���2������͏ߏ�� �%�4�U��j���r�����3��Ɵ؟��� �� �B�Q�r�5�����������4ѯ���� �ǿ=�_�nϏ�RϤ��Ϭ��ϥ�5� �� $�6���Z�|ϋ߬�o� �������ߥ�6�� /�A�S��wߙߨ���@�����������7(� :�L�^�p��������������1��8 E�W�i�{���;���� ��9 N���G �e tE�
� �  e���// %/7/g�V-�c�/+�/�d� ���/ ??&?8?J?\?R/d/ v.g:�?�;�?�/�/^? O*O<ONO`OrOh?z? �?�?�?�O�O�?�?~O 8_J_\_n_�_�_�O�Op�O�O�O�_ `F @� +e�/9o_Ywa�Uo�o�o�_ zj{o�o�o�o I[%/As�w ����!�?��'� i�{�E�O�a���Տ���\
Yo*���_MO�DE  e@�S �e��_�ZA�Uo~�П��	��� �CWORK_{ADP�
+��ȡ/R  er g���Q�_INTVA�LP���[�R_O�PTION�� �[��V_DAT�A_GRP 2�,�XpDPP�� ����C�1�g�U� ��y���������ӿ	� ��-��Q�?�u�cυ� �ϙ��Ͻ������� '�)�;�q�_ߕ߃߹� ����������7�%� [�I��m������ ������!��E�3�U� {�i������������� ����A/eS� w�����W���$SAF_DO_PULS;�X��A�Z�1!CAN_T�IMO�!U��BR� �(�C�(��f0/������Ē����S  �����//��7/I/[/m//�/���C,"2�$��)�d�$�!�&�@��\
??.?*��)�/ �ߠC4�_ 3b  Tf�W?�?�?��?�9T D�� �?�? OO$O6OHOZO lO~O�O�O�O�O�O�O��O_�����%_X_j_'Y+a��Q_;�o*����p(]
�t� ��Di�� -�� ,"���Q��y�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv���� �����*�<�N� `�r���������̏-��T?����+�=�O� a�s���ԏ�%��ß՟ �����/�A�S�X���-�0R2�S�U�]�� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� ߏ�ߪ߼�������� �(�:寧^�p��� ���������Y����� ,".�@�R�d�v����� ����������	' 9K]o���� ����#5G Yk}��������X�$_�3/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c?�q:0/z?�?�6������?�=	12345678�R_ !B�P
�8. �PO)O;OMO _OqO�O�O�O�A//�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ m�O$o6oHoZolo~o �o�o�o�o�o�o�op 2DoBHU }������� ��1�C�U�g�y���<��k;�j��ӏ ���	��-�?�Q�c� u���������ϟ��
iD���%�7�I�[� m��������ǯٯ� ���!�3�E�oi�{� ������ÿտ���� �/�A�S�e�wωϛ� Z�����������+� =�O�a�s߅ߗߩ߻� �����߰��'�9�K� ]�o��������������#�5�G�$ @d�v�[��������)"Cz  A��*   �(2`�4A��A!��0Ě22b�I[m����0/��� 8���!3E Wi{����� ��////�S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�?��?�?�?�$SCR�_GRP 1�(�ӈ�(ӑ �@t; �
 �1� 	 �3 AB	D���"M�7GJO8OqO���� nBD�` �D��C�GnK��R-2000i�B/165F 5_67890. �D�X. R2D7 ��@B#
1234��EAFnA� CV�1B&�3�1�DnAJBATY	ER��_�_�_�_�_�\���H��0�TG �2&o5O6o\ono=FM/
Io�oEo�o���o���h,P�Tn�t�� �AB���B��ffB�33B��  +v�5wAA��G  @
 _uAy@�@o  ?��w�rH-p�JzAF@ F�`�r�=GC�  ��� � �D�/�h�S���w�7q�_q�r������ʏ܄B���0��T�?�x� c�u�����ҟ����� ��*��CZOH�m���A  j���
�q@�p>��F��=G��߯-p���W\NCa�5�B$A�G�1Z��o��e �Y�
  {�����º��׸�\��Ŀ P�(!��'�9�K��1EL_D�EFAULT  �XT���
 _�MIPOWERFL  ��zw���WFDOl�� w�^�RVENT 1���`�u���L!DU�M_EIPM�����j!AF_IN�Ek��B$!FT$��>��b�!"o��� �Q߮�!RPC_MAIN����������VIS��ߕ	���F�!TMP9�PU=���d5����!
PMON_�PROXY����e ����Y����f��*��!RDM_SR�V+���g�v�!�R!T����he���!%
��M����i���!RLSYNC�5	8��Z!gROS�ρ�4Iަ!
CE[�MT'COM���k��{!	�CONS���l�>u�b9�/ A��w���� /�@///+/�/O/�a/Q�RVICE_�KL ?%�� �(%SVCPR#G1�/:�%2??"� 3+?0?� 4S?X?"� 5{?�?� 6�?�?� 7�?�?� TO<	9O K�$��HO�! �/pO�!?�O�!E?�O �!m?�O�!�?_�!�? 8_�!�?`_�!O�_�! 5O�_1^O�_1�O o 1�O(o1�OPo1�O xo1&_�o1N_�o1 v_�o1�_1�_@ B1�_�/�"� �/� � �1�����@� +�d�O����������� �͏��*��<�`� K���o�����̟��� ��&��J�5�n�Y� ��}���ȯ���ׯ� ��4��X�j�U���y� ����ֿ������0���Tϖz_DEV ����MC�:\���n�O�UT`�h��j�REC 1ŭuh���w h�	 \� ������<�'�`�n�
 ��u��XЃٛ� �߿߭���������� )�+�=�s�a���� ���������%�'� 9�o�Q���������� ����#G5k Y{������ �C1gy[ �������/ -//Q/?/u/c/�/�/ �/�/�/�/�/?)?? M?;?q?�?e?�?�?�? �?�?�?�?%O{�O[O IOOmO�O�O�O�O�O �O�O�O3_!_W_E_{_ �_o_�_�_�_�_�_�_ �_/oo?oeoSo�owo �o�o�o�o�o�o+ ;aO�gy� �����'�9�� ]�K�m�o�������ۏ �Ϗ���5�#�Y�G� i���q�����ß�ן ���1�C�%�g�U����y�������寽�V 1��� (ӯ&����TOP10 1���
 =�,�v������@�YPE��l�H�ELL_CFG ��{�h�Y� � n��B�RSR��/�h�Sό�w� �ϛ��Ͽ���
���.���R�=�v߈ߚ��/  ��%����P�ߨ�����b���L����װ�2b��d����϶HK 1�ݻ 
��� ������������� +�=�f�a�s�����������b�϶OMM ��ݿβFTOV_ENB���ƺ�OW_REG_U�I=ͲIMWAI�T:��mOUTr^�o	TIM^w���VAL~>p_UNIT9�vƹLCW TRY^�Ƶ��MON_�ALIAS ?e	�he:CXj |����R��� /�%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?�/i?{?�?�? J?�?�?�?�?O�?/O AOSOeOwO"O�O�O�O �O�O�O__+_=_O_ �Os_�_�_�_T_�_�_ �_oo�_9oKo]ooo �o,o�o�o�o�o�o�o #5G�oX}� ��^����� �C�U�g�y���6��� ��ӏ������-�?� Q���u���������h� ����)�ԟM�_� q�����@���˯ݯ� �� �%�7�I�[��� ������ǿr����� !�3�޿W�i�{ύϟ� J��������Ϥ��/� A�S�e�߉ߛ߭߿� ��|�����+�=��� a�s���B������ �����'�9�K�]�o� ��������������� #5G��k}� �L������1CUgy$�$�SMON_DEF�PRO ����� �*SYSTE�M*  ȏRECALL ?}�� ( �}$c�opy mc:d�iocfgsv.�io md:=>�portuc:8944�/)/;/M/�}.�frs:o�rderfil.�dat virt:\temp\���/�/�/�/]!&b&*.dv/�&�/?,?>?�Q-
xyzrate 61 �/�/�?�?�?�?Y%b7�+z? �?O/OAOT*1b/t(?mpback�/�O��O�O�O }(�db� *wO�H�O_._l@_S+,xbD:\�O�lP�K_�_�_�_W'-bUaj_|_ �_!o3o EoXOjO�O_�o�o�o �O�O�O�o/AT_ f_�_�_����_�_ uo�+�=�Poboto �o������͏�o{� �'�9�K�^���� ����ɟ�m� ���#� 5�G�Z�l�������� ů؏������1�C� V�h�����������ԟ �w�
��-�?�R�d� v����ϫϽ�Я�}� ��)�;�M�`�󿄿 �ߧ߹���޿o��� %�7�I�\�n����� ���������ϐ�!�3� E�X����ߎߟ����� ����y��/AT� f���������� �+=P�b��� ��������q /'/9/K/^p��/ �/�/�/�w/ �/#? 5?G?Z�/~?�?�? �?��{?/O1OCO�V(/�$:manu�tention.;tp�%emp�,O �O�O�OZ/l/�/O!_ 3_E_�/�/�/_�_�_��_�G�$SNPX�_ASG 1������Q�� P 0 '�%R[1]@g1.1�_i?��C%oDo'ohoKo]o�o �o�o�o�o�o�o�o. 8dG�k}� �������N� 1�X���g�������ޏ ������8��-�n� Q�x�����ȟ������ ��4��X�;�M��� q���į���˯ݯ� �(�T�7�x�[�m��� �����ǿ����>� !�H�t�WϘ�{ύ��� �������(���^� A�hߔ�w߸ߛ߭��� ����$��H�+�=�~� a���������� ���D�'�h�K�]��� ��������������. 8dG�k}� �����N 1X�g���� ��/�8//-/n/ Q/x/�/�/�/�/�/�/ �/?4??X?;?M?�? q?�?�?�?�?�?�?O O(OTO7OxO[OmO�O��O�O�O�D�TPAR�AM ��U��Q �	��JP�YTYP�XOFT�_KB_CFG � &S�U?TPIN_SIM  �[�4V�_�_�_7P�PR�VQSTP_DS�Bn^4R�_"X�@S�R �qY �� & �_/o&P�<VTHI_CHA�NGE  &T�\WOaGRPN�UMOV djOP_ON_ERRYh�ZY�aPTN |qUc`AKbRING_PRy`��n�@VDTsa �1�Ya`  	 8W"X0BTf x������� ��,�>�P�b�t��� ������Ώ����� (�:�a�^�p������� ��ʟܟ� �'�$�6� H�Z�l�~�������Ư ����� �2�D�V� h�z�������¿Կ� ��
��.�@�R�y�v� �ϚϬϾ�������� �?�<�N�`�r߄ߖ� �ߺ��������&� 8�J�\�n������ ���������"�4�F� X�j������������� ����0WTf x������� ,>Pbt�������?SVP�RG_COUNT�OV��a^U"EN�B�o	%M3#|eA/U�PD 1�kT  
�&R�/�/�/ �/�/�/�/??,?>? g?b?t?�?�?�?�?�? �?�?OO?O:OLO^O �O�O�O�O�O�O�O�O __$_6___Z_l_~_ �_�_�_�_�_�_�_o 7o2oDoVoozo�o�o �o�o�o�o
. WRdv���� ����/�*�<�N� w�r���������̏ޏ ���&�O�J�\�n� ��������ߟڟ����'�"�4� +YSDE�BUG y �K�d�a)l�SP_PAS�S%B?~�LOoG �x%c#�K�G�T�  ��]!K�
MC:\x��Z���_MPC���x%,�>�x!�\� �x!�SAV �b��Ф�G���SV_�TEM_T�IME 1�x)�
�(K��K���g"�T1SVGUNS�s %'a%�	�A�SK_OPTIO�N x%]!'!)�_�DI��4/E�BCC�FG �л�� 1���ψ�`��� ���������3��W� B�{ߍ�x߱ߜ����� �������S�>�w� b������������&�	�8�
�k�}� ��Z�����������c� ;���#I7m[ ������ �3!WE{i� ������// -///A/w/](H��/�/ �/�/�/]/?�/?9? '?]?o?�?O?�?�?�? �?�?�?�?�?OGO5O kOYO�O}O�O�O�O�O �O_�O1__U_C_e_ g_y_�_�_�_�/�_�_ o-o?o�_coQoso�o �o�o�o�o�o�o) M;]_q�� ������#�I� 7�m�[��������ŏ Ǐُ���3��_K�]� {������ß��ӟ�� ��/�A��e�S��� w���������ѯ��� +��O�=�s�a����� ��Ϳ���߿��%� '�9�o�]ϓ�I��Ͻ� ������}�#��3�Y� G�}ߏߡ�o��߳��� �������1�g�U� ��y���������	� ��-��Q�?�u�c��� ������������ ;M_���q�� ����%I 7m[}��� ��/�3/!/C/i/ W/�/{/�/�/�/�/�/ �/�//??S?	k?}? �?�?�?=?�?�?�?O O=OOOaO/O�OsO�O �O�O�O�O�O�O'__ K_9_o_]_�_�_�_�_ �_�_�_o�_5o#oEo GoYo�o}o�oi?�o�o �o�oC1Sy�g��v�p�$TB�CSG_GRP �2Շu��  �q 
 ?�  ��� ��@�*�<�v�`���謋�r�s��|d�0ہ?�q	 �HD)̪�&f1f�����B\�r��!��333?���8!�#��L�͇�L������C���ϖ��CAःC4����Ř@��  ����Ř���HA���@�p������¯���� �
�կ�5�R�a�7��p  ,	V�3.00�r	rw2d7a�	*��@���r��k���(�p7�� 㰵��  
�����M�&�-ÿqJCFG هuc�q�-��W����-ς�� �Ϩ϶ʐp������ � ��$��H�3�l�W�i� �ߍ��߱�������� �D�/�h�S��w�� �������
���.�� R�d��r�`o�����=� ���������� D /hz��Y�� ����q�A� QSe����� �/�/=/+/a/O/ �/s/�/�/�/�/�/? �/'??K?9?o?]?? �?�?�?�?�?�?�oO )O�?IOkOYO�O}O�O �O�O�O�O__1_�O A_C_U_�_y_�_�_�_ �_�_	o�_-oo=o?o Qo�ouo�o�o�o�o�o �o)M;q_ �������� �7�%�[�I�k���;O ����͏w������ !�W�E�{�i�����ß ՟�������-�S� e�w�1�������ѯ�� �����)�+�=�s� a���������߿Ϳ� ��9�'�]�Kρ�o� �ϓϥ���������#� 5�ߏM�_��ߡߏ� �߳����������C� U�g�%�w������ ����	����?�-�c� Q�s������������� ��)_M� q������ %I7m[} ��A���/�3/ !/C/i/W/�/{/�/�/ �/�/�/?�//??S? A?c?�?�?�?g?y?�? �?O�?+OOOO=O_O �OsO�O�O�O�O�O�O ___K_9_o_]_�_ �_�_�_�_�_�_o�_ 5o#oYoko/�o�o/ Qo�o�o�o�o/ UCy��[m� ����-�?�Q�� u�c�������Ϗ��� ���;�)�K�q�_� ��������ݟ˟�� �7�%�[�I��m��� ����ٯǯ��wo�o'� 9���W�i�����ÿ ���տ��/�A��� e�S�u�wωϿ����� �ϯ���=�+�a�O� q�s߅߻ߩ������ ��'��7�]�K��o� ������������#� �G�5�k�Y�����K� ����������1 ACU�y��� ��	�-Q;�  w{ �{�{�$TBJ�OP_GRP 2��C� _ ?�{	�ڮܵ�K�� `�pp� ���� � �< { @w�	 �D)�+%�C2
C랔�{�G"333O!>'���K/! LY p$/<��d+!? !p$�B`  A�A$�����'+/=/O%O"��/�*<+�~-C_  B�{@!�/?�/�/F'p%�%p={���5<ҙ*"P!p!�Cz!0�$�?��;C�6���C�p��.�?K��%p ;��:CA�ৃ"P$C�C4 �?VO�?�?m(�Oj;(A��=�/JhAH�0 �YO�OiO{O_+^ff=f?U<:f�/F ! �0?B�@f_x_+_�_�Y �_�_�_�_o�_�_!o ;o%o3oao�omo'o�o@�o�o�o�o"�D�{��  �G%	V3�.00�r2d7�*mp�v{��w GO ޛ~d� G�0G��� G�| G��: G�� G��� G�t G��2 G�� G��� G�l G��* G�� H�S�rFj` �~�� F�q � G�X G/� G�G8 G^� G�v G�ĺs��4 G�� G��� G�\ G�� =p =#�
"|8(1Cq�j�k�j}�{��?�X�����ESTPA�R�po��HR�րABLE 1ݒ���{���� (��v�������zT���	��
����T�{��������RDI�����!�3�E�W�i�єO ٟ�����+�=��	Sן� �����"� 4�F�X�j�|������� Ŀֿ�����0�B� TϚ֠گ	���~��� ����`�r�����������{�NUM  VC� �� �̐�_CFGG �d��!@��IMEBF_TT�܁ս逦�VER�ʓ������R 1=ߵ 8x{�v� F��   ��%�7�I�[�m�� ������������� !�3�E���i�{�����`����������_b̐�/ �  �k����T��>6���9��I���/ �LTA�_�6���Lu�6���Bx��� 7q����/ 
��E:��);^���g]o � �R�ƙs/� Vdà��/c W����
��/ [X�s!%�	/���_^����@��ӀMI_CWHAN�� �� �#�DBGLVL�����ҁ� ETHER_AD ?��� ��������/?ˈރ ROUT��!ƃ�!54S?&<SN�MASK�(���!255.�5Ys�?�?��?YsӀOOLOF/S_DI�pM%�)�ORQCTRL ���ɖ���1NT  OUOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�\O�_�_�_Ѓ�PE_DETAI��(�:PGL_CONFIG �d��tф�/cel�l/$CID$/grp1�_FoXojo|o�oD��?�o�o�o �o�o7I[m � ����� ���E�W�i�{��� ��.�ÏՏ����� ��A�S�e�w�����*� <�џ�����+���}��a�s���������)ѽ_�­����*� <�N�`�r��������� ̿޿���&�8�J� \�nπ�Ϥ϶����� ���ύ�"�4�F�X�j� |�ߠ߲��������� ��0�B�T�f�x�� ������������� ,�>�P�b�t�����'� ����������: L^p��#����� $`�E�User Vi�ew 4oXjI�}�1234567890��������@ c/��;2 q=/O/J�s/�/�/�/@�/�/=�//C3�/ !?3?b/W?i?{?�?�?�?�/�/<4�?OO F?;OMO_OqO�O�O�?�?<5�O�O�O*O_ 1_C_U_g_y_�O�O<6�_�_�__oo'o@9oKo]o�_�_<7eo �o�o�_�o�o/Apo�o<8I�� �o�����%�T�F� �ECameraFx��� �����ҏ�����E��9�K����x��� ������ҟ�`�+/� '���K�]�o������� �ɯۯ�8��#�5� G�Y�k�2�pu`�?�� ÿ������/�A� ��e�wω�Կ�Ͽ��� �����~����?M�_� �σߕߧ߹�����T� ��%�p�I�[�m�� ���ߐ��O����:� �1�C�U�g�y��ߝ� ���������	- ?��_����� �����9K ]������� R���o!/3/rW/i/ {/�/�/�/(�/�/�/ D/?/?A?S?e?w?� ����?�??�?OO )O;OMO�/qO�O�O�? �O�O�O�O__�?��9!_Z_l_�O�_�_�_ �_�_�_aOo o2o}_ Vohozo�o�o�o'_qt	a�0�o�o	Ho- ?Qcu��_�� ����)�;�M��o�l1Y������ɏ ۏ����#��G�Y� k���������şן�`��l2��/�A���e� w���������6���� �R�+�=�O�a�s������l3��˿ݿ�� �%�7�I�[�үϑ� ������������!����l4-�g�y߸ϝ� ����������n��-� ?��c�u�����4��l5����T�9� K�]�o�����
���� ��&���#5GY���l6e����� ��/��Se w�������<lz  w	+/ =/O/a/s/�/�/�/�/x�/�/�+   / 	/'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco��,  
s (  �� ( 	  so�o�o�o�o�o�o %'9o]��t�}j: �K �� ��D�V�h�z� ����u�ȏڏ�3� �"�4�F�X�j����� ������֟����� 0�w�T�f�x������� ��ү���=�O�,�>� P���t���������ο ����]�:�L�^� pςϔ�ۿ������#�  ��$�6�H�Zߡϳ� �ߢߴ����������  �2�y�V�h�z��ߞ� ����������?��.� @���d�v��������� ����_�<N `r������� %&8J\� �������� /"/i{X/j/|/� �/�/�/�/�/�/A/? 0?B?�/f?x?�?�?�? �??�?�?OO?,O>O�PObOtO�O�?�p@ A�B�O�O�O�C�G�`����O_&_8_ J_\_n_�_�_�_�_�_ �_�]_o o2oDoVo hozo�o�o�o�o�o�o �_
.@Rdv �������o� �*�<�N�`�r����� ����̏ޏ���&� 8�J�\�n��������� ȟڟ����"�4�F� X�j�|�������į֯ �����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφϠ�Ϫϼ����I(A� �O�$TPG�L_OUTPUT� ��1�1 ���,�>�P� b�t߆ߘߪ߼����� ����(�:�L�^�p������������  2345678901���� %�7�I�Q��2��x��� ��������j���,>P��}Z�� ���bt $ 6HZ�h��� ��p�/ /2/D/ V/� /�/�/�/�/�/ �/~/�/?.?@?R?d? �/r?�?�?�?�?�?z? �?O*O<ONO`OrO
O �O�O�O�O�O�O�O�O &_8_J_\_n___�_ �_�_�_�_�_�_o4o FoXojo|oo�o�o�o �o�o�o�o��}��0@BTfx��}@��������( 	 ����*��N�<� r�`�������̏���� ޏ��8�&�H�n�\� ��������ڟȟ�����4�"�X���OFF_LIM#���џ���t�Nw_SVx�  �����P_MON �َ���������STRTCHK ��Պ�-��VTCOMPAT���)���VWVAR �뿭"�N��� � � d���Ң��_DEFPRO�G %�%M�ANUTENTI�����ة_DISP�LAY#��IN�ST_MSK  �� кINU�SER�ִLCK�(��QUICKM�E��Nϔ�SCRE�k��*�tpscִ(����Ɋ����_��ST���R�ACE_CFG ���L�Ϡ	惴
?����HNL 2�L��S� y�?�Q�c�u߇ߙ��߽�����ITEM� 2�+� �%y$�  =<�xB�T�\�  !b�j�v�&���� 4����j�����i� ��������@�0�B� T�n�x�����Hn� ���,�P� "4�@���d ���L�p� K/�f/��/�/ /�/ $/v/�/Z/?~/*?P? b?�/n?�/�/?�?2? �?OOz?:O�?�?�? FO^O�?�O�O.O�ORO dO-_�OH_�Ol_~_�O �___�_<_�_`_o 2o�_�_�_�_�_�_jo o�o�o�o\o�o�o �o�ot��� 4FX�*��N�`� �l���Ï�ޏB� ��x�*����w�ҏ ������ȟڟ>��b� t��� ���V�|���� ���(�:���֯p�0� B���N�ʯܯ�� ��� $����Z��~���Y����S�����^��g  ��^� �����
 ��������d�R_GRP �1���� 	 @��L�^�H�~� lߢߐ��ߴޠ���߀�����%��I�4�?�  d�v�`��� ������������8� &�\�J���n����������	,��� )�S�CB 2�z� O�L^p������d�X_SCREEN 1�7��
 �}ipn�l/gen.htm�<N`r��&�Panel� setup�}�������/"/ ��Z/l/~/�/�/ �/+/�/O/�/? ?2? D?V?�/�/�?�?�?�? �?�?]?�?�?.O@ORO dOvO�O�?�O#O�O�O �O__*_�O�O`_r_ �_�_�_�_1___U_o o&o8oJo\o�_�o�_ �o�o�o�o�o�ouo��UALRM_MS�G ?7���� _zQc��� ������6�)��Z�M�~�2uSEV � @}��0rEFt��zϭ���A��_   B���� ��7��%�7�I�[�m� �������ǟ՗��1��Ƌ ?�4�����A��*SYST�EM*&�V8.1�079 G�1/3�0/2013 �A 7��5�"�U�I_MENHIS�_T   8 �$q�T_HEA�D��}�ENTR�Y ��$DU�MMY2  ڜ�3��  j�OU�SEt���$A�CTION��$�BUTTˤROW�͢COLUṂT�IME��$RE�SERVED���j�PANEDAT�t� � $P�AGEURL �}$FRA�)$HELP�{PA'�TER1+��<���H���H�4F�5�F�6F�7F�8+�I�NB�VA ���	�S'TAT*���1r���޸� j�US�RVIEWt� �<Ġn�U!��N�FIG��FOCU�S��PRIM!�m������TRIPL�*�m�UNDO_�t�t�  $�4�ENB��$W�ARNJų���_I�NFOt�y��_�PROG %$TASK_I���t�OSIDX��R���`�TOOL�t� 4 $X&��$����Z��ߡ�$P��R�°�N�U�9`�U&�t���������E��`�OsFF��u� D{�z��O?� 1���)�Q���GUN_�WIDTH  y��K�_SUB��o  
`�RT��t�t�	��$D�ܒ��ORN��RA�UX��T��ENAyB-���VCCM���� 
$VI�Sʠ_TYPɳCv(�RA��PORTФ��A�C���N(�%�$EX��_��$���_F�P��P� A���a�LU �$O�UTPUT_BMr�
���MR_�>��h ���<�+�DRIV����SET_VTC����BUG_COD~ɴMY_UBYȴ6�	����ʠE��,�ࢡ:�f�x�O�HAN�DEY��E�8pUL8X�P��AL_����GD_SPACI9N���RGT�������������U�RE$����U��w�������  ��R�G��PNT���R\���� dġXr��FLA���	T�A�XS���SW��_)A��y���S��O��BA��zy�	$E��UE���y�Ҁ��+HK�� �
зMAXvER��MwEAN�	WOR���z��MRCV��� ��ORG9pT_C&P )�
REF���- �i ��яN��b b1��_RC���� 8���M���M�ր��� �P�űG]�����$GROU�P����:&�� ���2p C�REǰw��$��Ab"N!HK��S�ULT���CO�VE����a NT6��%���&���&ձ�#m L6��%F��%����'ձ���9��0 &z#PA�u� z#CACHO�LOV*4@1��E9����C_LIMmIf3FRn8TDn8N�$HO��=�.0�COM������OB�O�8(� �!$IN�_VP�����2_S�Z3�#�56�#�51�2���8R��:TKQ��8o0�8WA5MP�BJFAIo0G��?0ADrIU�IMRyE $�B_SIZ/$�PM��ND� P�A�SYNBUFP�V�RTD�E�D�A�3O?LE_2D_��EmW�PC��TUq��@0Q� �EECCU��VEM��)54Ro6� ��$��� C�KLASv�	�V�LEXE5G���� �z!O�FLD6d�DE�CFI�@�W�� �W��;�s� a(����"R_ǠB�� ��_��L�#����Q�� hPP �1��!��K�$V��$=�E�!}ХC�U%$"A7
,�@PSKt4M:&�^e  ��TRb�Ut� $p TI�T-��A0=�OP�ɤ�VSHIF:�`��|!#�����URO�d _R �@�+tH�C=u��L� ^�p�o0���qi �ҏssTI�!�tSCO'r�sC����S¨�Sw S£vS°wS¾x���0�Ꞣ��s�ED���nw�  SM7��A���$ADJ,�`K��UA_{"u�qA��g}�LIN.Ӿ���ZABC������
!ZMwPCF��  C�d�J���LN�`p�a��I��� ��x�1� ��CMCM��}C�3CART_6���Pa $	JT�N�D�1Z�k�d�p��p����UXW����UXE�񞖙�_���u���������ɖ��ZP5��r��������Y��Dc� �y�2v/�IGH����h?(p ��|�$  � �d,7ۀ$Bm KK�]a�_�b�#u�RVn0F8��cOVC��O�@D��$�`��Ǳǡ
��Iݣ�5D�TRA�CEJ�Va��SP�HER�� ! a,p 1�G�Y��$��DEFx�?%����c��^�(%��x���t� ����ѿ������� *�O�:�s�^ϗϢ�T��IN��  c�ԢϦ�_T`H��1 �c�ހ(��� ��(/S�OFT͡/GEN���K?curre�nt=menup�age,153,�1��T�f�xߊ߀�9 �.�936A��� ������#�5�G�Y� k�}���������� �����1�C�U�g�y� �������������	 ��?Qcu�� (����'��ѶSew� ������// +/�O/a/s/�/�/�/ 8/J/�/�/??'?9? �/]?o?�?�?�?�?F? �?�?�?O#O5O�?�? kO}O�O�O�O�OTO�O �O__1_C_.@y_ �_�_�_�_�_�O�_	o o-o?oQo�_uo�o�o �o�o�o�opo) ;M_�o���� ��l��%�7�I� [�m��������Ǐُ �z��!�3�E�W�i� T_f_����ß՟��� ���/�A�S�e�w�� ������ѯ������ +�=�O�a�s������ ��Ϳ߿�ϒ�'�9� K�]�oρϓ�"Ϸ��� ������ߠ�5�G�Y� k�}ߏ�z��������� ����"�C�U�g�y� ���,�>�������	� �-���Q�c�u����� ��:�������) ����_q���� H��%7��[m��������$UI_PAN�EDATA 1�����  	�}��/ /2/D/V/h/ ) j/�/�$��/�/�/�/ ??z/7??[?m?T? �?x?�?�?�?�?�?O��?3OEO,OiOvI� ���B�/�O�O�O �O�O _SO$_�/6_Z_ l_~_�_�_�__�_�_ �_�_o2ooVo=ozo �oso�o�o�o�o�o
}L+v�H_M_q ����o�>_�� �%�7�I��m��f� ����Ǐُ�����!� �E�W�>�{�b����� $6�����/�A� ��e����������ѯ ���\�� �=�$�a� s�Z���~���Ϳ��� ؿ�'��KϾ�П�� �ϥϷ�����.���� ��5�G�Y�k�}ߏ��� �ߚ����������1� C�*�g�N������ ����X�j�(�-�?�Q� c�u����������� ��)��M_F �j����� �%7[B� ������/!/ tE/��i/{/�/�/�/ �/�/</�/�/??A? S?:?w?^?�?�?�?�? �?�?O�?+O��aO sO�O�O�O�OO�O�O d/_'_9_K_]_o_�O �_z_�_�_�_�_�_o #o
oGo.oko}odo�o0�o�o8OJO}��o !3EWi)�o� U}������ {8��\�C�U���y� ����ڏ�ӏ���4��F�-�j�v�TCNK�$�UI_POSTY�PE  TE� 	 v��͟��QUICKM_EN  �����П��RESTOR�E 1TE  �]�G�A�S�w�mr����� ��ѯ㯆���+�=� O��s���������f� ȿڿ�^�'�9�K�]� o�ϓϥϷ������� ���#�5�G�Y��f� xߊ������������ ��1�C�U�g�y��� ��������ߚ��� ��:�c�u�������N� ��������;M _q�.����& �%7�[m ���X���x/!/ۗSCRE��?�u1�sc<�u2\$3�\$4\$5\$6\$7�\$8\!��USER�> C/U"T= ^#ksTf#�$4�$5�$6�$�7�$8�!��NDO_CFG ����`�a��PDATE� �)�N�oneޒ� _IN/FO 1�&Q0��0%'/l?x8Z?�?~? �?�?�?�?O�?+OO OOaODO�O�OzO�OԜ�>1OFFSET ��OS5�� __0_B_o_f_x_�_ �_�_�O�_�_�_o5o ,o>okoboto�o�[ ���m
�o�o�HUFR�AME  �d�6;1RTOL_A�BRT932rEN�B;,xGRP 1�	0���Cz  A��s�q�a������v��*z��U[x1J{MSK � ^uQ3LyNq�%I:%�o��ݒVC�CM_PAp �
<%~VSCAM1 *ߏ�焣����5��V��MRwr2��ҀI�?��	с��	ֆ��Z�1B��5�A�@�pp�pȣ� 	�o����������<������uA����T�Z� B���o�Z�s� ����۟����ܯǯ � �$��!�Z���;����{���ƿy������I�SIONTMOU4:p^�˅���"�,��,��@�q FRk:\�\0A\�� �� MC�T�LOGa�   oUD1T�EX�����' B@ �������ϙ������ � � =	 1- �n6  -��� t������, ֌�_�=����h����z�TR�AIN��$�4��� (��h��ݧ� ���������"�4�j� X�n�|�����﯆/LEXE<��1�1-80��MPHA�SE  &53�k���R 2�
 ��]�o��������a������  ���� $6*1l����������� ��s����������G	no�pqrs�tuvw Z�~��� ����./f</ n`/r/��/�/�/�/�//h$/?H/&? L?~/p?�?�?�?�?�? /? O2?$O6Oh?ZO�lO~O�O�OD�{u�3��? �OO__LO>_P_b_�t_�_D��D	��BH
�O�_�O�_ o4_&o8oJo\onoH��@~		�3�
�
��Æ�o�_ �o�oo&8J�|o�3�
�
ghijk�@ \��o��o�o����&�8�ƃ��SHI�FTMENU 1,>�c�<��%�ϖ�&���t���ӏ���� 	����?��(�N��� ^�p��������ʟܟ �;��$�q�H�Z����~�T��[�K��	VSFT1��~VSCAM�S�5ذ?��!�@`��G�  A�ٰ8*ٰٰ��p*�$����"�!����9�L�̦MEP �a�/� T�MO����zR�WAIT?DINEND � �|w���OK  O�ȵ��ԿS迻�TI]M����G�� 5�ǿX��8��8�%���RELE9�h�s�f��TM��s����?_ACTIV��1����_DATA 	[�2�%��h�,���RDISg�����$ZABC_GR�P 1۩I�,�qp�2p�t�ZMP?CF_G 1�v��I�0�������MP¨�۩/��'��8��'�s�8����0��_����?����� ���/����V�������`�[������@�������Ѕ������P_CYLIN�DER 2��� Н� ,(  *m~��j���� ��% gH�lSe�� ���-/��D/ +/h/O/��/�/��=�s2 ۧ4� �� �/<�~�3??W?e:h�/�?�7��1A�;�SPHERE 2!M�/�?R/�?O �?8O�/�?nO�O��O CO)O�O�O�O�OWO4_ F_�O�O|_�O�_�_�_��__�_oo��ZZ�� ���