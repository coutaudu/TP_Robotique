��   a�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����PASSNAM�E_T   0� $+ �$'WORD  �? LEVEL � $TI- OU�TT  &F/�� $SET�UPJPROGR�AMJINSTA�LLJY  ?$CURR_O��USER�NUM��STPS_LOkG_P N��$�eT�N�  6 �COUNT_DO�WN�$ENB�_PCMPWD �� DV�IN�!$C� CR=E�PARM:� =T:DIAG:)|�LVCHK!>FULLM0��YXT�CNTD��MENU�A�UTO,�FG_wDSP�RLS�� �$$CL(  ? ���!���	��	�VIRT�UA� /�$DC�S_COD@�|��%�  W6'�_S  $*�!$& t&�A91F"%!�N 
 $ !���-�/�/�/�/�/ ??,?:?P?^?t?�?��?�?�?�?�?��#SUP� �+�?�?�#�FO&OfO��  �L�A���O� � �� V�?[t&��j�� �B3O�O��G�O��/X.U.V