��   �A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����FSAC_LS�T_T   8� $CLNT_�NAME !�$IP_ADDR�ESSB $AC�CN _LVL � $APPP  _  �$8 AO ? ���z�����o VIRT�UALw�'DE�F\ � � �����ENA'BLE� �������LIST 1 ���  @!H������
 [.@�d��� ��/�3//W/*/ </�/`/�/�/�/�/�/ �/�/??S?&?8?J? �?n?�?�?�?�?�?O �?�?OO"OsOFO�OjO |O�O�O�O�O_�O�O 7__\_B_�_f_x_�_ �_�_�W