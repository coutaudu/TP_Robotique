��   j�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����DRYRUN_�T   � �$'ENB  �$NUM_POkRTA ESU@�$STATE }P TCOL_���PMPMCmGR�P_MASKZE�� OTIONNLOG_INFON�iAVcFLTR�_EMPTYd ?$PROD__ L ��ESTOP_D�SBLAPOW_�RECOVAOP�R�SAW_� G� %$INI�T	 &J_ � 4 $TY�PENFST_IcDX�@_ICI�  �MIX_�BG-1
_NsAMc MODc�_USd�IFY�_TI� gM�KR-  �$LINc  � �_SIZc�g� [. , �$USE_FL�C ���i�S�IMA�Q�QB�&'SCAN�AX�C+INC*I��_C7OUNrRO���O!_TMR_VA�g�h>� i �'` ��B���!�+WAR�$�mHp!k#N@CH���$$CLA�SS  ���� 1��5��50VIRTU� ?00'|/ >55���U����w8?0'1~5��%'1�?���?��?��O5I1Z; �O&O8OJO\OnO�O �O�O�O�O�O�O�O_`"_4_�?*W?>5{d1 ��Xt_�_�_  �1~0��_ k 1Z;G 4%B_�_��{1 �1�_%ooIo[o:oo �opo�o�o�o�o�o�o ! W6�1�S��Z=�9~0�� �r~1�tX{1>1~0�> ����*�<�N�`� r�����������~6�1 �q�1� ��$�6�H� Z�l�~�������Ɵ؟�$4v6�S�1Z9 �)�;�M� _�q���������˯ݯ ��Ό�4�F�X�j� |�������Ŀֿ��� ��0�B�T�f�xϊ� �Ϯ����������� %�>�P�b�t߆ߘߪ� ����������!�3� L�^�p������� ���� ��$�/�H�Z� l�~������������� �� 2=�Vhz �������
 .9Kdv�� �����//*/ </�6