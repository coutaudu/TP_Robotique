��  �\�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A9  �����ABSPOS_�GRP_T  �  $PAR�AM  �  �ALRM�_RECOV1�   $ALM�OENB��]OyNiI M_IF1� D $EN�ABLE k L�AST_^  �d�U�K}MA�X� $LDEB�UG@  
FPCOUPLED1� $[PP_P�ROCES0 Խ �1��UR�EQ1 � �$SOFT; T_�ID�TOTAL7_EQ� $,�NO/PS_SP�I_INDE���$DX�SCRE�EN_NAME ��SIGN�j��&PK_�FI� 	$T�HKY�PANE�7  	$DU_MMY12� ��3�4�GRG_�STR1 � �$TIT�$I��1&�$��$�$5&6&7*&8&9'0''@�%!'�%5'1?'U1I'1S'1]'2h"�GSBN_CFG�1  8 $�CNV_JNT_�* �DATA_C�MNT�!$FL�AGSL*CHE�CK��AT_C�ELLSETUP�  P� HO�ME_IO� }%:3MACROF2�REPRO8�DR�UNCD�i2SM�p5H UTOBAC�KU0 ��	DEVIC#T�Ih�$DFD��ST�0B 3$�INTERVAL��DISP_UNsIT��0_DO�6�ERR�9FR_F�a�INGRE5S�!Y0Q_�3t4�C_WA�4�12JO�FF_� N�3DEL_HLOG�2�jA��2?�1k@�?Q�� ���H X_�D�#	 d �$CARD_EX�IST�$FS?SB_TYPi� �CHKBD_SE��5AGN G� �$SLOT_N�UMZ�APREV�D�G �1_ED�IT1
 � *h1G=H0S?@f�%$EPY$�OPc iAEToE_OK�BUS�oP_CR�A$�4xJVAZ0LACIw�Y1�R�@k �1CO�MMEc@$D�V�QOk@:Y���$QL*OU/R , $�1V1AIB0~ OL#eR"2�CF�D X �$GR� � S!1�$MB_@NFLI�C�3\`
UIRE�s3��AOMqWI�TCHWcAX_NR.0S�=`_;G0� � 
$WARNM'@f��@� sLI? �aNST� �CORN��1FL{TR�eTRAT@0�T�` �0ACC��1�` |�rOR�I�P�CxkRTq0_sSF� �!CHG]I1 [ TT`�u3I*pTY��	RpK*2  x� �`� 1�B*H�DR�J* ��q2��v3�v4�v5�v6��v7�v8�v9� ���CO�$ <� Mo_oqh�s1<`�O_MOR./ t 0Ev�kNG� �0BA�  �Qt�Q}��r��@�!�v���P�0��XQpA0�f�`^P@/P�2� �p�JpC_R�bLq�@�J	rL	�$�JV�@�CD�`�m|gv�uMtP_}0sOF� �  @� �RO_����aIT<8C��NOM_�0�1���q3� ���$ !����|hP���mEX�`G�0� �0"�<�`�b
$TFR�J6 �D3��TO�3&@yU=0�� ��YH�2�T1m�E��� �e��f��f���0CPDBGDE���@$`PqU�3�f)����AX 1�dbET;AI�3BUF�F��|���! � ˧��`PI���P�L�MK�MX���[�F>L�SIMQS��wKEE��PAT�`��!� �����MC�U� �$}1JB8�`-�}1DEC㺋���ԓR� �7PCHNS_EMPvrG$GA�'��@_y�<q3�`1_FP͔x�;TCR�SPEubw�@q0�cg�S�!�� V�A0���!����JR!0��?SEGFRApv �r�R�T_LIN�C��PVF�r������Y��P���)B��وD ) \�}f�e	�"��	�ఀ.0�Z��Ql��SCIZCuх�d�To��A��ڭ�	�RSINF��p����?��������s���LItx�1���CRC�eFCCC �`��>�R��mRMAl�R��P� �$�D�d�c��C��j@T�A�����@��l���E�V���jF��_��Fw�N�� ��f��!��� 2���������1C��! ����h#RG�Ps�
qF��7b�g�D���2g�LEW(��s� �e�>�P��PqR�D� �&�pou2|��A6�NHANCI�$LG�`-��1�Pd��@�dB�aA?@l���~0R��z�jME��uAk��feRAs3jAZC���T�OEqFCT�q��`F�`m�g�̰�ADI;�  q�� l��`��`�`|��H�S=P�r��AMP��Ĥ�Y8C?�MACES����r�I�$�  *�I���CSX�a�!M�p	$JTpT��X�C_ N�@h�IMG_HEIGH�A��WID��h�VTtE��U�0F_A��8- �@EXP(�cN-%�CU���QU�1w $`TIT�19RISG1ꀿ��?DBPXWO���0= �0$SK���2�� DBT% TRN�@ !^�Q0TC�؅ `��DJ�4LAY_CAL�1iR� �'�'PL	3&@�0E�D���'�Q�'�QȘ"��!"�"1�PR� 
� �q��!g# T A$wqS$�љL@9$M?H_3Gp� %s?�4C�!9&�?�4ENE�ax�c'�?_3!0RE�`��2(H C�p �#$LC$$@@3�B� K��VOa s_D6G�ROS�b�cvh�D��AMCRIG7GEReFPAyS�>��ETURNcBo�MR_o�TU�`\)�2@EWM����cGN`��CBLA����EΑ�P��&$P� 9�'�@�QU�1C�D���0DO�����-DAS�3FGO_A7WAYCBMO���Q�m� CSC0EV}I>@ ) HJ`�1vRBw���SPI�hpJ�SP`wVI_CBY��|S�UHSL�r�*XP$��avVTgOFB�\�dFE=A�1v�SvTHS�+ �8��DO?��cnpMC%�d�P��)b�R����! `�,� $���J �c #fc ��faסߠebit�c�H�fa�"afWr��dNTV�fbV-pr��� ؃���g�s?�J�?�<�0��SAFE̕v�_SVq�EXCL�U�!����ONLd+�<sY�TktOT!!���HI_V5�PPLY_,�etw�]f�js_M8� $�VRFY_�#�O�� �v!1��s�b8Fc"�Q -�0� r~�_�:� vGaSG� .�
$���@�A����U�REV�-�$��UN�0xK�vU��턍��@��l�i�!Xq����rEFf`I�2/��$FN�X$��OT�@jS$DUMMY
1ׄ1ׄ�����M�PNIG20C L����4���A`a��DAY�e`AD�iT� ��؃5��EF( $���1�0ѧ��Y�_3� _RTRQ�ݑ2 D_�Ot@R�Q:���'���Y� 21����~�jT|�8�s�¡3 0��ؑ �	�גS�U�@]��"CAB¡4��x��$��$ID��CPW��ӕH�g�ViW�V_Ӑ��0�DI�AG�q¡5� '$$V�@a�T�ǃ� ��� ��
0	�R�25���VE� J�SW������(���~����2ZP~�OH���P�P���IRs!	�B ��7�����Aᇀ��BAS9q�z ���HiV���4����Cנ��RQDW�MS�9���A�������L�IFE� ����10��N��
�ɵi���
�h��^Ui�Cm7Q�N�@Y����FLA�Tj�OV6նHE<���UPPO��w	��� _6�� , �6 `�pCACHE-�m��Es�B~�SUFFIX��e`� ��@�R�؃6\ԁ�rMSW�7bKEYIMAG�C�TM%AH����A��I�NPU�?�!OC�VIEʠ�!8 �h�� L�d��c?�� 	�!"�9���$HOST� ! R�
0Z�0Z�G�Z�R�>Z�EMAIL\ E��� SBL��UL�G2:"҃�COU���T�T�0y�;' $��eSӐ4�;IT1cBUFǂaP�NTf j 5�B�ԂmTC�dA��s#��S#AV<��҅�EK@b2W�Ppm�PC�e�0�ˤ��_��"�`��OQTRBu�?P�pM�e����r��Z͓DYN)_�� <��DtU� ҀU���TR_IFS�W�O��A�!=0��/�Ӡ�#$@TIKYD#&��L�A����K���/�D�SP��/�PC��I�M<���sM�w�U`f�+�XE�p��IP�cd/���DC`��TH0Ȱ|�TLA��HS<��ABSCH���	F��s�dk�$���o�SCi�ʖ�1�!�!>6bFUI�DU��c�f�@PE���CD��	 ���W�R_NO�AUTO�!?��a$���:�PS��CC`�C�"s���q��� @H *�LI ���jU s@�c>
1<1<@G�<R�<��<79�8999��;E1�R1_1l1y1��1�1�1�2����GR`�Hl2�y2�2�2�2*�3�3E3R_U3l3y3�3�U3�3�4�sXTz�NaA <�� �� �]V �jU��7���FDRi�?BT ��	���ò�17òREMr��FQ̲OVMb�z�5A�9TROV�9�DTG�JMX#LI�N�98PJf�IND�2@ʲ
^H* s�$DG
�X+�@M`ɵr��D��@RIV�U�̲GEARb�IO��K�2ʴN$��HY�स_p�`�a̲Z_MsCM��ñ �F,�;URwC ,�Wq�?  �p?\0P��?0QEop28QD`�aCOԐO`�D��n�P1av�RqI�QTz�UP2�p3E G���TD��os��S0�HQ�W�U�zUB;AC��F TP���T�Ł)]qG�U%��8� t IFI�� �XP]`+��UPT̢.QQMR2�5G���1�s�2LIxaFc�7��O�O�OF��ʵ�2_��N��_������M�F�O�MDGCL�F�DGDYxL	DHQ�D5Ѷ�Oɴ'c�E�Hϐ�i T��FS��F�I PแxqL`
�s�$E�X_wq�xwq1��E�Zwq3�{5�v�GsRA�P�4J ���tSW%�Ot�DE�BUG�#���GRt0���UZBKUe �O1  ΰPO`0��CԐ�t��MS�`OO��^�SM�`EK�����0_E K S�|�P:��TERM��yL�����ORI`�M����SM_��P�҅�N�����T�AǉO��� �UP>�P� - ��2�K$���L$S�EG�%pELTO���$USED�NFI�<�Pt�� |��
�M$UFR�R���� 6�����`OT���pT���0��NST��PATx���OPTHJI� EH�s� �=�AR��I���8V��<�REL�r�SHFT =���ۘ7_SH:�MO�Ɔ� р��5�O�a�0O#VR��r�&�I��d5U� ^�AY��Q`
��ID�MhS�� q� ERVDx�7 &� h2������!`ӥ�!�`RCXQr�ASY1M"�r�=�WJP�h1�d@EhSב�����U�'�������ђ�P�����V�OR��ML@c��GRo��tQ�� �U���l���W�S�E�_R � h�QTOC6�:�Q��OPbm���*tv�e�1OA�RE���RT�r�O
�]⮒e�R��>����T�e$PWR�@IM0ũ�R_���S�]�w S�P$H�U�[�_ADDR�6H�r�G������vѷR�=p��8�T H�pS ` ���#���#��_���lSEkq�IF��HS� �sU $���_Dm0=���6+�PR��z�ð�TT��UTH7�V� (� OBJEC�a!(Q�Q$�6L�E��_�8�W�px7��AB__A�Գ��S��I�DBGLV���KRLp�HIT�E�BGD�LO����TEM���%B��g�SS�@7�HQW�C���X��\��INCPU�rVISIOR���Di����j��j�l �IO�LN��Y} �@C��$SL��$�INPUT_u��$0���P�@���S	Lp��Z������{IO@�F_AS]r[�P$L�P���QD-�.Uƀ)�T��� ���z�HY�7T�-���UOPZu\ `�r�6BBD�B@K���B�P90�����K�������J�6] �� �PNEV�JsOGk���DISBc�J7/�OF�$J8	7W IT�'97_LAB���) �QAPHI�`�Q(mDypJ7Jx��0�p_KEY�` �Kk��0\s^ �@��V��{6��CTR퓵FLA�G�rLGʴ_ ��9`y8���sLG_SIZ�ԧPXp,�FDI" Q�
��	� �Xp���9���<�2@SCH_H��R�� N�r`~�����p�q��1�`U�H����L#�DAU%EAP�k�ܴ3"�) GHݲk��BO}O�Rat B3��IT�3g$�`/�R{EC|*SCRN� �/�DI.�Sl�=pRGMb�0�,��'����"$���S���W�$��$'�JGM7MN3CHF�'�FN�6�K;7PRG99UF�G8W�G8FWDG8H]L~9STPG:VG8�`G8n G8RS�9Ho�c;$�CY��3&�'��p�'IUG�[4�'H���&� <�N2G+9�PP�ORG�:�%�3P/6O�C$�J8EX#�TU%I95Ii�#�B�# �C3�C70;11���AC��'1��!NO�FA�NA�6��`VAI�Q ��CL�a��DCS_HI	�NR��MR1OSX�aVTSIxWjX9SvX�(IGN"���481�  `UUDEVL���BU`��b� �_�T�B$EAM�[����3A��c� _���e�W�Q`*m@19e29e39aR$9_}Q��d ����`{�5���%��IDop�X�.�4�=a�&���fSTs�R4 Y�p1��`� c$E�fC �k��F��f�fXfo���e LL�B��pW�)� � �C����PЄ��"~�#_ f :�@�V����!�s|�C��g ���CLD�Ps���TRQLI�i � �y�tFLG �b�p�a�s=QD��w�=�LD�u�t�uORG �2�r���8����ҙt0�h � �	�u�5�t�uS��TD�p� s�!�����RCLMC��<�N�0��������MIН�gi d�yaRQ� =s�DSTB���`c ��!'�AX���� *�C�EXCESH�a��MO���j�P����q��Nџ�k���_A����A�S��pKʴl \�L��$MB>�L�Iw��REQUI�Rˢ
��O�DESBU`B��LSpM��m��4�Z������F��ND	!ǰ��n������DC�B$INeЫ!$�� ���P�N�b�C�PST��� o��LOCf|fRI&�|eEX��A��}a���ODA�Q�p
�$ON�RMF�@`��i�RrJ@\u����SU�P��qFX�IG}Gz! q �s�@Rs���RsFRtR��%�cιs�޸s��<ΐ<�DATAg*�EEq�E��T�N�R�r tN�MDK�I�x�)YƎPd��a�H�/�"dĸ�Ue�AN�SW�!d�a�Ad�D�&�);��󔀟�s -��CU"V���p�7�RR2��t���Z���A�� d�$CALI ��GtAQ
�2��RINP0��<$R�SW0�ʄH�y�ABC_�D_J2SE4��X��_J3s�
m�1S�P?�< �PmԔ�3P���������Jy���Մ�V_O�QIM<y���CSKP�z�H�:S�J<!��Q��3��3�)�$�_AZ����e�EL�Q���'NTE��"bu����7���%p_N��v@����a���䛒w��3DI{���DHc���:��x� $Vв�v�a$;1$Zb�N`b�����yH �$S v��TqACCEL�Q�U�ׁd�IRC��T�?�T�a�c$SPSc��rLn������s��z��BP{�P�ATHZ���p���3���f�_6a$� 䙂M`C��k�_MG�!$DD${�"$FW��=�`�@�p�k�5DE^PP�ABN��ROTSPEE:a��p)�:aDEF!�k�n��$USE_�SP��CO@SY� 6�- ��YN �A� ����{��MOU!N�GO� OL��INC��,�]D'�=<��(�ENCS�#�`���k�%���IN�b�I��>���)�VEx"Ӡ23_U�b�LOWL�Q I@���pi�D,@� ����Wpi��C���gMOS�PӔMOܰ�����PERCH  �OV� �1'|a <#�a����a2�m"� ,����P��A��%LT��З�ך�����&�TRKE$�bAYLOA���"�� 1���53-��`S�RTqI��K�`MOM�B�'���2����\
�03��9b5�DU�����S_BCKLSH_C��5&D ���°4d�:+�CLAL`���A0���5�CHK�p�eSRTY�@(��@�e$�r<�_�c$_UM��r=ICJC$SCLWDn� LMT��_L6���pE��|GEvM�@�K u@���E���Ц1
� L�Du(PCB!u(HYp�;�(@EC��]rXT\k�6CN_%�N�SD7V׃S�P� g(V���c|V�Q��{UXC!`HMSH�c%�6l $�{1{�2���U��f$PAGD;_PFE*3_�pd@6% �q3)dEJGxpy�c��OG*Wn2TORQU� ��# 9l ��"�o1l �b_WY5 4_@�e�e�eI�kI�kI�FE��a��Xx]�. VCZ�0!��"r1(~u�<2�/u�JRK(|mr`v��D�BL_SM7��Mΰ�_DL�GR�V�d�t�t�qH�_�S�s���zCOS�{/0�xLNop
�+u ������aH�6���a�uZ�&�qMY�����rTH�}��T�HET0�NK2a3�т��CBֆCB�C �h����d0	��	�ֆSB�'�N�GTS���C�� ,��S&��PS�6�`�E�$DU@И��
� G������]1Q�2�'$NE䗰I�(CH�2R���$��ŁAɅ�����u�x�qLPH�uВ�ВS'�C�6� C�E�ВT�m�W�t���EV�V	��,�V;�UVH�VV�Vd�Vr�V��V��H�-�3�P+��QJ�H�HV�Hd�UHr�H��H��O��O�O��*�O;�O�H�OV�Od�Or�O
��Ot�FВ��R�6��W��SPBALAgNCE���ALE>�H_ɅSP��'����6���E�PFULC����½���E���1u�LUTO_@=eTg1T2�V�2N�1 q�)�6���:1�������U1T� O{�c�`�INSEGq��R�EV���DIF��%��1v����1w�� OB���1�sg72�x`)�A�tLCHW3AR��AB�Qi5?$MECH����X�(FAX1P�Dp,�����x 
-⸋aO�|ROB% C�R�"o�!R��MS�K_��9�z P !�_� RV�����$1zR����ػ4����IN|��MTCOM_Cp>=�{   ��~v$NORE��������| 4�`GR�b�FLA�|�$XYZ_D�A�B`��DEBUb?� ��$�} ���$�COD�1 �o�>2�90$BUFINDX� ����MOR��~ H��W0e��6���5�4��J��&Q��@TA����g2G�� � $SIMUL'`�v�X#�#OBJ�E��ADJUS<1$ AY_I>az(DROUTG`>�W0n_FI=��T�`�	��I��Ф`�� ��в��%D� F�RI�3�T�5RO�g`�E�a� �OPsWOnp���,|�SYSBU⠙�$�SOP���1U<��PRUN��<PA��D;�s a_m �B1��ABc��@m IMAG�14�ฐP��IM���IN�pd�RGO�VRD�- oP0q�xP��L_	ЄQ��<BWPRBXP��>�AMC_ED��� �@N�M"�A�0�MY19�A��S�L����� x �$OVSL[�SDI� DEX@SR&OS$�!p"V�`m%Nw!�a�j� u#�'�(%"AQ�0$_SET�`���� @�`�"6�1RI�0
�&_��'�!��!���/ lP ���T�<`ATUS>~0$TRC��� ���/3BTM87"1I�Y#$4�A3 ��� D��EmV",2렁E��-1�� �0-1EXE30)A!�2�2f4b�#�� ��20UPI��1$�ИXNN�X7q#$q[9 �P�G�� � $SUB!16��!!1�#�JMPWAI�PPz#9ELOy@9���$RCVFAIGL_C��RP<AR�   �)�QjPATs��E���R_PL�#DBTqB<anRRPBWD~Ff�UMl`�DIGT�<ћ�
BDEFS}PH� � L���3��@_�@7�CUN!Ir]7�@�1R�0�r�p_L��P+1�C����k�e`�q� J�t���N��KET@R��`W�HPP�B��� hB ARSIZAEw�:� I�QS/ �OR�#FORMAT��DCO5 �Q~��EM%��T#SUX�� �"�BLI�B���  $��P_SWI���Eqp�@�@�AL_ � $H�A���B!��C���DY$E�1��,`C_�A� �� �@�d��(aJ3xr����TIA4�iu5�i6��MOM��@�c�c�c�c�c��BP@�AD�c�f�c�f�cPU
�NR�du�cu�b�!�R�� C$PIǖoe��od �tWu�sWu�sWu��v@m{ �r�[!P�j!{��$�6�SPEED��Gb�tQE�D�v�D QE�@� �v��x�A��AQESAM����Z�8�w[�QEMOV�򊔀���Л��������@1�䶄2��� ��`��d%`�H<Т�IN� %`>�����QB�2�x	�2�R�GAMM~�|��I�$GET����;D_d��
1�L�IBR�1GrIT�$HI�0_�;0��ǖ�E��ԘAΞ��LWɝ���3��[b.%�MTN+aC�E�����  $PGDCK�$�;_=� � ��$bph$a؅���c����f��)c �+$I� R"�D�����1rD��LE����!��[h�n`MSW�FLY��T�И���Pq�UR_SCR��3`�-�#S_SA�VE_D�~��3NO_`C�!�2`d~��� ojXv��qy��0�� ۻN���v�̀Ja`  <����љ��������x �v��|�x�6Û���1*tM2u� � ��YLQs��؇Pр��ɣ�Ǟc����W��w�����p��d���M��(�CL'؀(aC&"l�"&�q/!P�LMo��� � s$���$W~���NG�ya~�8d|� ?d|�Fd|�Md�@���P��c�%`X9POGc�$aZ��P@ �� pB ��ʣUv��ҿ������_a_�� |B oi~��i��c���c~��j����jE�@ ���U��U��\�tz`��P�Q�PM� �QU_� � 8�TPQCOU̡^ Q�TH��HO��c�H�YS�PES��b�U�EN�t��POd� �  ���"UN\40*� 
@O���� P���oE`�|}3GrROGRAG1
��2�4O����R��ސ�INFO�� ����� ����AO�I#� (R�SLEQ�vK�uK �����D>@����O������sƑE�N9U��AUT���COPY���0�j!
��M�N� �m�C�� �QRGADJʢᚓRX�R$P9P.�.W,P,`$�.�s&CEX�@cYC��1NSD�� � $A�LGOz���NYQ__FREQ��W=�0�v��T�#LA��pѫc=��uCRE�0̚#� IF�"��NA6c�%�_G�&3�(%���ELE-@ {�jbENAB���PEASI_!|� ��N"�q���&cBՀ��I ����qf�_`�&�"AB�!K`E���p9V��'BASUb�%౒���0���0$��!6��� X� �" 2� ����>62=7;QX�ޠR5i6�B�-P�F��RGRIDd�13CB�P�wTY`#N�OTO���@���_$!Z�2C$O� ������[@P�ORqC�3Cv�2SReV )	DFDI�P�T_�p#@5D��?G3�=I"P?G5=I6=I7*=I8!A�@F�������$VALU��#q�r$ �A���| [%�����3!n��PANp�vS0 1R�0�Qn�TOeP`�,��$SPW�I�1:TREGEN8ZMROc�X7�s�v���FI�T1R�#1B8Q_St��WMP�#Vѵq�U�q<!#GRTb�Q�Slì�ܯ SV_H�0DA8Y�P�PS_Y������So�ARY�2��+0CONFIG_SE_�PBn�d2���G�5� 4W�?�v�v[�6�PS~���{ @W�MC_Fl�|�a�L�~��SM����a�bNs�����c� ,R�F1L�Г���YN�`|UMf0C���9PU���LY�ᦛ�DELiA4pb�Y��ADY��� �QSKIPN�ŧ ľ���O��cNT��o1^pP_�� ��}w`��ҵ��w�Q�y �Q�yV@�zc@�zp@�z@}@�z�@�z�@�z9�qO�J2Rf���fbEX��T�C�n��C��0rC���q�R�DC֩ ���R 塘�M�ͅ����f�w�RGEA�R� ]�`�E�D��ڝ�ER�ar^�C~UM_C�~p�J2TH2N��~4� 1� t��EFI�1�� l�(�4�\#����TPE���DO�]� ����T���O3S���ՒP��~��&�2.��4�@F�X�j�|�����3.����ß՟������4.��.�@�R�d�v�����5.������ϯP�����6.��(�@:�L�^�p�����7.������ɿۿ�����8.��"�4�F�X�jϼ|ώ�SMSK��B#�
�'�bPD�5s��EMO& ���f`0�6�V4�IOT��I���P1�POW;ER�� 6�ppa����S ��e��$DSB� �!�T/pC� �RS2�32:ն� *�D?EVICEU�". |t�RPARITY�.!OPBITSF7LOW0`TR�� R+P���RCU��r �UXTASK�RINx�FAC��1"�і��CH���b�`_�sC����POMx�tbPGET_�@ �b� g0���P[��߸� !��$USAp�1���� O�`� ��'`���_ON�P����'WRK����D�P�~��FRIEND 1x $UF��#w��TOOL~�MYH��`t�LENGTHw_VT��FIRM`ȧ��U E�е�UFwINV ��RGI�MAIT�I�r��Xzq�� G2 �G1�1U���d+�0_y�|O_�� ����#� ����@�TCs��D��QG߀1#b`��`�� ���bo
�.%�S0#�R� �������XS ��v0L�T�H�0��&����)$IW�0�EDRpLOCK6'Aqwp�Q�Ui�Q$�20����4�.�:�1F�5�2*8�2�38�3F�� �G��!�����S��R�SV�P��VVV@��� �`b`��� b��so:�|+e $p�qP]P�! ��S���U����A9@�'P!R�P�&��SS�q� ��q���2� 0��0�20�haV#�������E U�{r
��S^��� �c!RA,Q{2$P`N��`�BHAn�L��rw2/THIC.� pap�C��TFEREN�1t5I�@H.�w1I08��3��K0G1�(�4����9�r��6_JMFGPR�`}q�b��C� <q� *R �}r�C �-F{� ���ҢA  2� ��Sx����	d' �$��Du��Ep�C$Pn4�CDSP�F�JOG�P�p`_P�q:�O�1Fu��� L�7KEP��IR�A�D2]`MUAP&�!E�%P�4�S`�@��R�PG:VBRK�`�5�0n0I�� A aR�clR�Br A�R<�C�@BSOC�FJ�uN�UD#`Y15�q�$SVDE_�OP9dFSPD_WOVR�a<pC�`L�R�COR�W��N��b�VF�1�V�@OV�ECSFjP`c�F3f��!�CHKh��"LC�H2rFuRECOV(�T���@W"pM�P�eF�@RO8�Q�@_h0�a0 @���VE�R�p��OFS��CN@��WD�Q�d�Q�QX��U�PTR,� Ѿ#@E_FDOVMOB_CMb�	pB�@�BLs"�B+rs!�$V@�	��� ucbG,w?XAM=SpZ mu�b�_MCpE�ހOӹ`OT$CA�@ހDhR�pHBK��6�q�IO8��upсPPA�z��y��u�u�pҹbDVC_DB ��C��1��D��b�![�1c��s[�3c��`ă�U��@�QUK�@O�CAB�@7��� �ch� fx
�OzpUX�6?SUBCPUr2�@SQ��sUt��*#��3#Ut���Q$HW�_C��D@pH�A�.c0�$UNIT�uTo�h�ATTR�I-P|��@CYCL�ycNECA��SF�LTR_2_FI`�4�خ����1LP�K��0�0_SCTvF�_h�F_r�����FqS��Mrm�CHAQ���<�Lr:�;�RSD��`�҅Q�3s1p�_T�jxPRO��s0�E%M��_�`iST)�:!� )�C!��DI����4RAILAC4Q��Mz@LO�P���T7t� ���!���s+PRE�S�10��C7���	�cFUN9C�R�"RIN� s�02�Ġ:�/�RAK��� �pc�p�tc�W3AR�3�pBL|y��A��������DA`sPd�θ����LD�� �P���o1m��!���TI�"�xac0$���RIA���AF
�P�Aä`GŶ8[S�ʓMOIs�v�DF_��Jc��C@L�MOsFA��HRD]Y�ORG��H]��v2�ְ��MULS�E��-S�L!��J��ZJ�Rg	kFAN?_ALMLV,���WRN�HARD�`в��� ��n�2$?SHADOW`�0���AMU_�`�6A�U� R.�F�TO_SBR9��յ@��h��9�B���MPINFBa0~������5��8p�`|A�  d��$!�$�� �xBbA}@�� ��2SEG���C�P%�AR�@���U201躰�?UAXE�GROB��FW��fQ_t�SS�YrP_�hP��S��W�RI��8�*!G�SCTR�E��gP�PEj��K@A�oҽ B���a���!�P�pOT�O��K@�`ARY�n3+�䡘�UA�AFI�HP�C$LINK(��~1K�/!_��a�@��!r�XYZt:�}�5��OFF�`RJ�r�f�/�B�@�/����a��3���F�I����:1�R�T/��D_J�AIB�RW�`e����S�TB!d��YC��.VDU�b\?���TUR�XÈ�9��X���pAFL0 g`ǃ2� ����y8�R�a 1�K@%K�@M�4?�9���8�"��cORQ���Ai���3H� EP�0��Э!`-S�ATrOV	E|�2M��1�Ӗ �Ӗ�IГO�� j��E4��H��1} �@�d��1�}�%0��%��AER�Am��	��E��1@�]$A!c0��[���7�ձ҆ձAX�cIBձ�� Q�L�%���)���)�� �*���*�P�*���*� �*�*1H��&���) \0�)\0�)\0�)\0�) \09\09\0/9\0?9�\1P9DEBU@��$;�Gӯ� A�bn�ABէ�q�Qv[@Ġ�r
Bl�7!CEb�OG� OG��OG��OG�QOG�� OG�OGM�^ G��.��LAB��A<��I�GRO��A@��pB_��D&���S������F,QB(U��4VAND� ��R$��w�U!��qW �q��v�XƱ��X��v�NT'��:>��SERVE�P�� $��g�Axa!�PPO�b��p%��Q�S_MRA��/ d ԰T�`xd�ERREsC�TY.���I�pV��#2a'TOQ�$�Lc�$���Ee�T�C� � px ,P�d��_V1^2�!�d���d�2�k2�f�QW�� �8@@�Q�s$W���f�TldV����$`���w��"jeOCƱ���  kCoOUNT�� �Q�HELL_CFG��� 5 B�_BAScRSR� AB��#�i�S�j��cp1�U%bq2��z3�z4�z5�z6ʆz7�z8�wVqROaO���pݐu�NL���dAB�S͠dpAC-K,FINpT�4���e���.��_PUXՓC��OU�SP���guܡDr�v��чTPFWD_KAR7aLc aRE�T��PG�ܱ��QUEm���}���A�c�I�/CCs�s�ڣ?�v�at�SE�MR�	�b���<�.PT�Y%�SO�!DDI�1����Cс�'u�_T9M�P"�NRQb�s��Eߐ C$KEY?SWITCHڣ���D�ڄHE��BEAiT����E5�LE6b�����U��F����S~I�DO_HOME��OO�REF]PR���"����2�CԐO��`qaO�P3@�&��IOCM_�YA�@wHK�� D<p�o�RESUbς�M����ooFOR�Cs�ʳ ibDsO}M6� � @
DT=Â�U��P4�1֦��4�3֦4�ibN�PX_ASKr� �0qpADD{�Z��$SIZa$VqA2P�u��TIP�)�۠A���`` _�����]�S�C�yC2`y�FRIF���pS��˩�i�NFpe�
�dp�� xx SIObTE�P��SGLѱTY� &�����C��ҰSTM�T��P!���BW<}ӴSHOWř���SV�����; �	aA00vTT� ߠ\��\��\���\�U5Z�6Z�7Z�8Z�9Z�AZ�W�\�ʠ\� �A]���\���_�O0تf�1s�1��1��1���1��1��1��1���1��1��1��1
�1�1�G���f� ���؀ɉ��ؚ�Q ��P��� ����2��2��U2��2�2�2٨V��f�3s�3��3���3��3��3��3���3��3��3��3���3�3�3�4���4f�4s�4��4���4��4��4��4���4��4��4��4���4�4�4�5���5f�5s�5��5���5��5��5��5���5��5��5��5���5�5�5�6���6f�6s�6��6���6��6��6��6���6��6��6��6���6�6�6�7���7f�7s�7��7���7��7��7��7���7��7��7��7��7�7�7�v@qVP��UPDJ�G� �`� {r
�P�YSLOKr� � #�i�f���� S �4R@U5;�Ԏ�pR@8F�!ID�_Le�h5HIc:I���PLE_b��4��$	��&SA�b�� h`�0E_BL�CK���2���8D_CPU�9$��9�c3��?�4�"P]�R ��|`
PWp�q -FALA��S�aKC\AUDRUN�ErAJD rAUD���E�AJD�AUD_ �TBC�CJ��X -$�ALEN��D��@?��RA��R� W$PI���F1�A�42WM�p]��C��.�ID� 9jQ&\TOR�@�>[D�a0S��LAC�EB�0R�@c0R6`_�MA	�MV�U]W�QT#CV�\�Q]WTn��Z �U�ZСKT�a�U]S�a�JA�
t$Mdg�JH��D�LU9a]U�A�2A�<��`RaKS"PJKefVK�wa�wa�3icJ0�d{cJJv�cJJ�cAAL{cP�`�c�`�f4�e5�B�QN1�\�`�[�P.T%L'P_��>�
@p�@�Is� `�0GR�OUN0�g�B��N�FLICa�=pRE�QUIRE
�EB�UJ��AfY��P2��X��@]v�A�G��{ \m�APPRipiCT��P
��EN�x�CLO��yS_M�����yLU
�AL�7� �7�MC�R�P��B�_MG���C�F��0$�␉P%�BRK#�NOLS�%�2�Rc�_LI%�i�S��Jr�e�P�diP�c�iP�ciP�ciP�ciP6��߱��8B�\��B�t�� fr�B�A� ��A�PATH 
�#��#��H�N�xpm�dPCN�CAt��i��r�IN�BUCh-P1y�C�PUM��!YPl���l1E�@����@���`o�PAYL�OAa�J2L� R'_ANx��LG@���ߙ��$�R_F2�LSHR��%�LO��x�)���7���ACRL_�v�i�r�הr�BHA0�R$H$�ޗ�FLEX�s��@J�E� : �O�F]Pȧߤ�O�A]P�O�O\F1ߡ-�A��_)_;_M___q_q�E {_�_�_�_�_�_�_�_ oH�e�g$cedU�w� ,o>oPoޡWjT��F�Xl�bce����ne� �zo�o�o�`�e�e�e@�e�o�o�oyrJ!t� � -?Q���� ATZ�eq`EMLȰ *�lxJS���spJEP�CTR,r�U�TNv�F(�]wHAND_VB�q��M0�� $���F2$��sb�<2SW�A6r�v�� '$$M��R>���@O������厂�Ao0 ܐ�n1$��A.�10
@�AN�A]�/�/��0�@�DN�D]�P=�G]@��STB���O���N`�DYt@�p$�� 7��}��ߡ�:�ޗ eg�����d�P���� ��Å̅Յޅ��Ӓu� �ത���<�q�ASYMM��	fpM�ۤ�h�:�m�_SHrw���{�@�蛟����џ�J���������g�_V�I����s	 V_�UNI/�$?�'�J fe6"d6":�:$Q�G$ k&Z�`m���|����%�������1q�pH�H@�rݙ��!ENL��
�DI]���O4q q� !s� O�
>�I!A��Q�819@��3F3�08��p;A�1�o � ��ME�����a2�"HT� P�Tq��8��1pt �p��8�1�9T�q� $DUMM�Y1G�$PS_fX�RF�0$�6m!ALA#pYP����2�3$GLB_T��5E�01�@��Y�'1� X�p]w��ST��spSBR�M�M21_VbT�$SV_ER�O�Wp_CwCCL3@_BA�ɰO;2� GL  E�W$q� 4+p�1+$Y�Z�W�C[`$$���Ab0���"�@]U�E� ��N�@�v0E$GIi�}$�A �@�C�@$q�� L+p�Fr}$yFrWNEAR���N_�FLY��TAN9C_��AJOG?���� ���$JO�INT�!q��EMS;ET$q�  �I3T�ʱ��SM�U��$q����MOU��?��spLOCK_F�O9���0BGLV�\�GL�XTEST�_XM�p�QEMPĈP��b1B�P$cUS~1�@� 2�sp��C@a�b���P@a��aACEpSa` $�KAR�M3TP�DRA�@~duQVE�C�fyPIU@a��EaHE�PTOOL�!��cV �RE�`I�S3��d6ÁU�ASCH�PS���aO[�ԑ3�42�PSI��r  @$RAIL_BOXE�!�spROBOd?��aAHOWWAR�0q�0�aROLM �2Vu���dgr��p�Td�a��_�DOU�R� H R^cI�2���P$PIPfN���br�ag�@a�p�C��OH0 �{ D�pGLOBA� 6��P���3@�r�8�SYS�ADR�7�� �0TCH�� o� ,��EN�"*1A�Q_�Dp��Ѿ��PVWVAd1� � �`�B5PREV_RTq�$EDIT��V/SHWR��KFԀ���A�Ds0
���HEAD�� �����KE�A�0C�PSPD�JMP�_�L 5��R��#4U��e�I`S7�C}�NE�`8�s�T'ICK!�+M�ѵ�F�HNAA� @p�pc���$�_GP���v&@STYj��aL�O3A�CF������ �t 
��Gv�%$ԕ��D=K@S�!�$,!� x1E50FP��SQUx`�B��TERC�0��;TS��� �&AW@@�ר���x��aT�O�0��3c�IZD�AE�1PROC�2Ѣ1�pPU#!�_DO�QRo�XS�PK 6A�XI �zsEaUR �ɳ8�7p��.����Y_�`@�ETA�P�RT����F�
t��R���l  ����ꔵ�榹� ��� ���0�ڵR�ڵ b�ڵr��͟��*� �
��s��C)�k�}���t�SC�@ � h�@D1S��a�0SP20�AT`��⡠�o�~�2ADDRES�c=B��SHIF��7`�_2CH7�*�I�:@X��TXSCR�EE����T�INA�CPk��D�rPB��C@� T U�z@Ţ8�yAV@���p7���Լ�RRO; �fP7����W4�AUE�$4� �� Y��0S��A8�RSM���U�NEXk� 6"�� S_�CB�%2�E�`�%�B�C�R�� 1-�t�UE{��,2�B\��ѠGMT~ L�!��f@O�V�$$�CLA<� ������0�@����V�IRTU� ����A�BS����1 ��� < ��9�K�]�o� ���������������� #5GYk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?^=���AXL�������+�  �p4IN�y?�1o4��_EXEr�8�0�6_UP���1#���LARM�"�OVoP��2l4L�M_P���d^?BOTO fOxO�J0O�O�O�O�O�M, 
6�_j6�NGTOL  �#�	 A   �L_^[�PPLICf��?��0�P�Handl�ingTool ��U 
V8.1�0P/11  ~S-C�(
ya�SW�RՠԄ�Q
F0�Q�U����ՠ
1232��TOh��X��Z��`��7DC�1�P\�SNone�  EL@T�FRA_ 4��YWbl�PpQ��TI�V�5�S�3�cUTEO�� A�4�9P1�GAPON��n���`OUPL�p1I� �`&tg9�`UB� 1K) ��0x0|0|�����s�1�s���� ��Uvt�H_ur�zHTTHKY���cu� ���#�}�G�Y�k� ��������ŏ׏��� ��y�C�U�g����� ������ӟ���	�� u�?�Q�c��������� ��ϯ����q�;� M�_�}���������˿ ݿ���m�7�I�[� y�ϑϣϵ������� ���i�3�E�W�u�{� �ߟ߱���������� e�/�A�S�q�w��� ����������a�+� =�O�m�s��������� ������]'9K io������ ��Y#5Gek��|BuTO6P�o�cDO_CLEAN�o|@t#NM  ;[_Q/c/u/�/�/4�_DSPDRYRL/?uHI�`/-@@/ ??+?=?O?a?s?�?��?�?�?�?�?<xMA�XrP����g�1X���Q�b�Q�bPLU�GG�`��c�ePRUC� B- �+�/��?WBO\B�/@tSEGF�`K�O�G�A-/ ?/__+_=_O_�O�ALAP�/�N�s�_�_ �_�_�_�_o!o3oEo�Woio{o�cTOTA�LFHI�cUSENU�@�k ��o��BpRG_STRI�NG 1�k
��M�`S}j�
q_ITEM1v  n}m6HZ l~������ �� �2�D�V�h�z����I/O S�IGNALu�Tryout M�odeuInp�̀Simulat{edqOutތOVERR� � = 100rIn cycl҅�qProg A�bor�qȄS�tatuss	H�eartbeat�wMH Fauyl\�e�Alero� ��������ß՟���8��/� �{ �(2���������ȯ گ����"�4�F�X��j�|�������ĿF�WOR�@{��p�ֿ$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D�8V�h�z�PO{P� ��ˉ���������� �/�A�S�e�w��� �������������DEV��D��1�k� }��������������� 1CUgy�����PALT \����"4F Xj|����� ��//0/B/T/�GRI@{�! f/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?z/�`R\�0A �/
OXOjO|O�O�O�O �O�O�O�O__0_B_�T_f_x_�_�_OPREG��PHO�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
.�@���$ARG_���D ?	�����q� � 	$��	+[�x]�w����y�vpSBN_CON?FIG �{ց�Ղ�qCII_SAVE  ����q�rvpTCEL�LSETUP ��z%  OME�_IO����%M�OV_H9�L�R�R�EP3L��pvUTOoBACK$��}�FRA:\��[ ���V�'�`:��W� {� �� �x �]>�P�}�t��������������� )�;��UΟg�y����� ����L����	��-� ?�Q�ܯu��������� ϿZ����)�;�M�_�>A��dωϛϭ�p�����ϲ�INI� ��T�u��MESSAG����p>�ODE_D>���͆9�OF�H߶�PA�US��!��{ ((O�r�߲ۜ� ����������*�,� >�t�b������{�~��TSK  ��x��Ϲ�UPDT?���d5�U�XSCRDCFG 1�v_������|��������� �����e�0BT fx����������rs��G�ROUN)�i�UU�P_NAf��{	���R_ED�1�
L�� 
 �%�-BCKEDTA-Cz���[��P�����Z�r��xW��r/  ��_%A2h/y�F/�/<"��t %�/�/C/U/�/y/a#34?�/�?�/�.]?�? ?!?�?E?a#4 Op? MO�?�.)O�O�?�?�OOa#5�O<O_`O�.��O`_�O�OO_�Oa#6 �__�_,_�.�_,os_�_o�_a#7do�_�o �_�.�o�o?oQo�ouoBa#80�}h�-�Y��Aa#9�lI�4��-%���`����a!CRg/ �o�&��m�Z������I�׏U�NO_D�ELasGE_U�NUSE_qLA�L_OUT ���>#tWD_AB�OR��T�IT_R_RTN׀l��NONS���.�1�CE_RIA�_I)�5�y�FFF���.���_PARAMGPw 1�����?
��.��Cp�  O��Q��Q���Q��Q��Q��Q���Q��Q��Q��Q���Q��Q��  D���I�p����y�����둴� D���Ѱ��"Ѱ*j��1Ѱ9��@�.�?�y�HE��ON�FIG#���G_P_RI 1���� �$��S�e�wωϛϭ�ܿ���CHK��1�5� ,5��� %�7�I�[�m�ߑߣ� �����������!�3�E���OF��찫t�CO_MORGR/P 2֬ h����� 	 �������������̣������q?����p�`�R:Kh�:��Pa�������a�A-��������.
��
��r�@����.��`MCPDB�c����9)c?pmidbgN��� �:��s�t����p�����U�^ �^ ����-���t��0�v�����Egf��"Ff�/��/� mc:,/T/k?DEF "(��)@ cebuf.tx��/�
a/}��_MC��u F԰ d�%�#���-��!5Cz  �BH�B���B��H'B�`C��B�r-C�Z���D3�6C�G�C���D@OC���kD�w�Z=E���E�OE���\E�dE���	F��	?G�����%4����<	j��4~*j�������A3x���C\Q�D�Di�D@Z>N@� DE�D�  F��E�oF�`/R�> �JBE�L@Gb��FO��\G�L��:� � >�33 �9���;  n��;F�5Y�E��; Aa��=L��<#ׄ�2i�E�O/�"R�SMOFST �.���)T1��DoE �� ��Y
�Aj�;��B�O��O�.TESTy"._v�R��g��_%6CC4�@���� A!�A62��;0Bl�;0�C(@@c��j�:�d�
�QI_����]�QT��FPROG %,���o�UT_IܑZ@䖏���dKEY_TBL�  6��
A� �	
��� !"#�$%&'()*+�,-./0123�456789:;�<=>?@ABC�y GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾�����q���͓��������������������������������������������������?��������z`�L|��kp�z`ݐSTyA"��T_AUT���Oe��V>�IND�T_ENB+���ROQI�;�T2��t�a��n���XCˣ 2��j��8
SONY XC-56�_�	B�u��@�����  ( А{��HR50
Ȓ��+�7=�O�ACff[��o��ß �� ���՟�0��T�f� A�����w���ү������f,TRL|`LE�T��� w�T_�SCREEN �,�kcsc���U��MMENU� 1u < *�o�������S ǿ�&����\�3�E� ��i�{ϡ��ϱ���� ����F��/�Uߎ�e� w��ߛ߭�������	� B��+�x�O�a��� ���������,��� b�9�K�q��������� ��������%^5 G�k}���� ��H1~U g������� 2/	//A/z/Q/c/�/��)k�_MANUAyLÏF�DBCOe��RIG4�5�DBN_UMLIM��:��d�UY`DBPXW�ORK 1 fk��_[?m??�?�?�]D�BTB_)� !��_�Q�PK4�!_A�WAY�#:�GC�P �R=|P�6_A!L0-��2�"Y6���P�(_DBG 1"ZY�I�,�K?�O��SrO�O�8_Md�I�)PL@+`�CONT�IM3���T���F?I
�eTCMOT�NEND�oSDRECORD 1(fk� ��O�SG�O�Qm_�[B�_�_�_ �_xX�_o_4o�_Xo jo|oo)o�o!o�oEo �o0�oT�ox �o����A�e ��>�P�b�t���� ���+�������� :���E�͏�������� '�ܟK�՟o�$�6�H��Z�ɟ~�i�w����@e�served f�or Tool  �����m�"���X���@mmy $0E=0u� #33Y�������ƿ�������@	�! TP Key2 (ABOR�@ $�6�HϷ�l�ۿe���k Pq�5u�9 گ ����X���ώ�C��A�t Release)q�8u�E�|ߎ�����JTOLERE�NC DB�IB@L���� CSS_D�EVICE 1)>�9  �6� �)�;�M�_�q�������C��LS 1*���������!�3��E�W�����PARA/M +`Ii�����_CFG ,�`Ki�dMC:�\��L%04d.'CSVh�� c��i�YA��CH z� ��Oi�Q���'��2�!~l@0�J�PѦ�RC_OU/T -�;m@k�~��SGN .�5�?R��\�1�6-MAR-22? 15:01��?1z� 4�4:45���� Tnu��-)i�*�o���Im��P�uG��=��VERSI�ON �
�V3.1.j�� E�FLOGIC 1�/�; 	�(�@0����PROG_ENB!OFR�WULS�G �6��_ACC6(A��.C�7#WRST�JN�@�&?R�#DE�MO,(A0E{!IN�I� 0�:�5?1 �v&OPT_SL �?	�&�"
 	�R575i�� 7U4�)6�(7�'5j�
2182�$�6?�>�$TO  �-@t�?�V� DEXd'�d?U�3PATHw A�
A\�?��?O�KIAG_G�RP 25���� �	 E� � F,D FAD�`QC��@IC@��nO�LkA��ЗO�NCe�ECl^OCk�I$C��C�� B�m�I�f362 67�89012345��B�'  �cP�A���A�=q�A�A�33�A�z�A���A��RA���;A�P���JPj!@\@p	 GQ���A�������B4�L��D�(j!
R�P�{A�P��P؜P�P�G��Aď\A��A�Q�*?_Q_cTP�*�б)�^�PϸPU�P� P��P��P���A�ffA�P#P�_�_�_�_o��X_�PZ@`U�PO��
AJPDP>*$P8P2@`,�lWo�io{o�o�]`��A�[�PV�PPPK
=AE�A?P�8��A2�P+ׁ
�o�o�o�X���`�$PLpxPq�Pj$Pc P\Q�;ATPL��bt ����TC@R�Q3a�aKq�p^M=�G��z�>8Q솅^M8���b��7�Ŭ���^M@ʏ\ʆ��p�օE@[PAh�	 �C@<�C�<��t�=�P=�hs=���P�^M;��
.�<#�8�[ �?+���C�  <(��U� 4Ƃ�̝�r����~���@
"?fE6���8���� ��9�k��0�ʟ@�f��H�����~�?Tzᐾ�;�ʥ^M�{��G��^NcQ����^Nx`��7��C��O
�@��CkJ=C���Ck�^M�m����|��ఱ`K
�׿%�ED � E�� ��D+�	�C��O7�j!�8�?6д�����9b�V���6в�eWZ�2����b�����DkC��耚���#Ϡ����{������I ACT__CONFI��6������eg�� ASTBF_TTSd'
)B�C#t��U���MAU^ \/��MSW��7���_P��OCVIEW�i�8��	 �� �����*�<�N�I ��~��������g� ��� �2�D�V���z� ������������u�
 .@Rd���� ����q* <N`r��� ���/&/8/J/X\/n/��RC��9�5v�!
/|.�/�/�/�/��/#??G?[�SBL�_FAULT �:�*��a1GPMS�K�7t7�0T"A �;ٵ���M�C: �C�O�:|#P ��OO1OCOUOgOyO �O�O�O�O�O�O�O	_8_-_L� ����1ORECP�?�:
�3 �_���?�_�_�_�_o o,o>oPoboto�o�o��o�o�o�o�oI_��U�MP_OPTIO1NK�m>qTR��L�:q9;uPMEJ�.�Y_TEM�ï��3BK��p��ytUNI��MՏq���YN_BRK �<��y8EMGDI_STA�u���q��uNC�s1=�� C��o'��|,d�_ m��������Ǐُ� ���!�3�E�W�i�{� ������ß՟|+��� ���[�&�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���2� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� ���*�<�N�`�r� ������������ �&�8�J�\�n����� ������������" 4FXj|��� ����0B Tfx������ ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? ��?�?�?�?�? OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_�?f_�_�_�_�_ �_�_�_
oo.o@oRo dovo�o�o�o�o�o�o �o*<r_`r �������� �&�8�J�\�n����� ����ȏڏ����"� XF�X�j�|������� ğ֟�����0�B� T�f�x���������ү ���,��,�>�P�b� t���������ο�� ��(�:�L�^�pς� �Ϧϸ������ �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/��/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO �/�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6olOFolo~o�o�o �o�o�o�o�o 2 DVhz���� ���
��Ro@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟ޟ�� 8�&�8�J�\�n����� ����ȯگ����"� 4�F�X�j�|������� Ŀֿ����0�B� T�f�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������ ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������� �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?��?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ x?f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o L_&L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���2 �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ���*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶���������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x��������� ������,�>�P�b� t��������������� (:L^p� ������  $6HZl~�� �����/ /2/ D/V/�f/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�?��?I�$ENETMODE 1>r%��  _   4@4@�<E7OIH@RROR�_PROG %�#J%�LH�OLFdETABLE  #K�|/�O�O�OJRR�SEV_NUM �2B  ��-A)PdA_AUTO_ENB  PE�+CaD_NO>Q �?#KEA(R  �*��P��P��P��P4P+�P�_�_�_ZT�HIS%SLA+@S[_�ALM 1@#K� �LD�\�@+ �_;oMo_oqo�o�o�_�_R`P  #K�QFB�j@TCP_�VER !#J!��O�o$EXTLO�G_REQ�V�QY,sSIZ5'tSkTKRyoU�)r�TOL  LAD�z�R�A 't_BWD�`�pHV�qDww_DI�q Ar%�STDDLAKB�vS�TEP��@�pO�P_DOtbAFD�R_GRP 1B#INQd 	�or�F@�c��[��w���#/[��7u���� �����c����ɍc�C�?B���NB�!B�z�A�O�B��N΍B���B�l��BMӯA�f��A�YA|��΍ɏ?�*�c��N���r�����  A��8A��>煖���D@
 �JN$&�֑Β�Cv�b��ׄEݐ�F,D :�D�`�E���)�D  Ew�� b�D+�m�{C�(�C��N���B�ƈ��΍@UUU��UU��ۯ&�~8��� E�@����΍OHcGP{)�K��6�/Jk�΍?�R���:G:�z�9{󨂆�΍�����t<���n�LA��������KFEATUROE Cr%�pJA�Handl�ingTool �� svde�English �Dictiona�ry��
! �4D St�a�rd�  ffs~��AA Vis� Master���� R597�nalog I/O(ǿ  90 HS�g�le Shift�(�R6417�ut�o Softwa�re Update  4 RR���matic Baockupe�49����ground �EditI�  o�adiCam�era[�F_�4�t���nrRndImܸ��duc��om�m@�calib �UI�� ERm�C�on��@�onit{or��ct\j3��tr�Relia�bt���PCVL�Data Ac�qu=�:���.sv�k�iagnosx��X���cflxk�ocument;�GeweE���'�Ok��ual Chec�k Safety�%� g H5��h�anced Usf��Fr���PC���xt. DIO �5�fi�� def�.��end��ErrD�L�������בs-����rV��� �p��41m�FCT�N Menu��v�`���H55��FT�P InF�fac�v�  J�JG���pB�k Excz��g�� Par��T��Proxy �Sv��  j61�6�igh-Sp�e��Ski� 6�.fd㰎��mm�unic��ons������urm�F�_�? R67\����connect �2��04��Inc�r��str�z�F�CB��KAREL Cmd. L���ua��J�Uc�Ru�n-Ti��Env�#�"
c�P�el� +��s��S/W���  �L?icense�Ӳ����$�Book(S�yE�m)��! t�oMACROs,��/O3�{���IF��H���
 �81 ��Mech/Stop��t:�z�o T "j�Mi�rw� ����Mix��xX����orch���odu�witch�(���o:҉�. �d -��Optm� R7*����fil��Pick��X�g� OAD~�ulti-T�������v
EPCM funT��z�90#ow�Re3giE��  d����PH�t F* D�/�[Y�Num S{el6  ry��|y�� Adju�����k�w�  p=r�tatuR*�GNDI��ٵ�r���RDM Robo}t�scove�N*�Rem4 �n�� ,���	#Serv�o� ��?SNP�X b��(�rt <�w�Libr���Gpbo��w�� EN{   m� W o��tm�ssag �Pv��!z�[s in VC&,Ӧ��`q ���(TP�"�/I�� )��� M�ILIB=fxt�p� P FirmĖ�)�d���n�Ac�c����e�71TX���L��� eln <I0� �����e\mc�1rqu>u�imulaC���_ te.f�1u� �Pa���Ma��T���^Ѡ&��ev.��Ѧ�USB po�o @�iP�a�� ���,@nexceSpt��# n�� ��\@�����n0VCb!�r���:hk�1�<�j4<�{+�4<�S?P CSUI��l���IXC�&ro�H�x�� 
�W�eb Pl���9!7��QC!�Nl21R����ԩ�D��3%F� �i�gXGrid!play o�gX� ���L� �iRnIV�MRe  e� -�2000iB/1�65��rAsci�i���1�� 5 ;(K�UUpl��񷤣35�s!��!t� ;rc��Cyct����]ori��5%FR�L��amY*�HM�I Dev�� (Y!����PC��-@o >#asswo&�2
�49\��64MB DRA�!	�l2�b�FRO�kY�7�rcN�visD���5c����ell[�L�H5M4�sh*q�"�0�C|c�^�2@Eu��pX�6JDEutyt�s���VIct�� .���� ��sp 2���aV�B by �
 ��	 B"X�q i3t2���T1>�K%�.10�OL�`S�upB�Rc�O'PT ��njNS �b9S�B�cro��cx	#{%�T mjp��x='�a�puest*��SS�`e�tex�{� ���$LimipYb�Sp����1��0P���gJ�n�Virt��	#���M�dpn�8��h51�>CVIS� IR�pvC�JDIRCA�Lv>D�+�IC:�;0x ��phi�cD�hо�Abui4�l�� F�!�PMM�p�� !fwlowh1f.sk�OSFILE A�r" u�co gt�p��BMON��IgX c�җ!m T��N@PTTB:��i��R805� ��J����
��⊔j��^�m����"PAL{T:�`clud����AIW�- Wa�it/Y�ea�� �tk��TP�bDO�ES NOT R�ESTO �60L{in��markЎ�useJ�z ��c��  Synchr�@�z���DSUPP�R��PRG INW AR�A ��Ag���OVC_VAL�UE�OBLEM� ��V��TMi�TMW��G���ab��A MOTION��STRUCT �l��BRAKE ABNORMx�� ��g�$FMS�_GRV0ISMA�TCH=uu�Z�MA�ST HANG �UP 37m�MU�LTI WIN/�LOCB���SER�VO��AG GA�R*�
�GRID �DETECT B�UA���!0�����T�RANSLAY�OF UTX���F DB/s�DO� PULSE@E�NCCAMERA�ǁ�c�`REMA?RK FOR�� �w�L�0\h���E�XPANDED POS>���%'�|���SCREEl��AY CRUSH� �P!�OTN5�60����fԡ�ND��SYRUNNIp��Ɛ�USR���F TOLp�NC�E ��vK�FSE���Ŧ ���S-1�44 A��ARTؾ�
p�FA_� CPMO-073�w�AUIs�0��mp�l����ڢ�ps�ᇡ�����R��sydem�ַ��A~��snosv.�Ј���޷�i���gA �S���HQ��a_cUmC�-PH�T���!  ORsPAd&;6�`�PR��r[qdp�(Co��Y�P,�" �1�ҷ���G���ҷ�g�R5c56�ִ���ic��`e�|��G��tg���2�G���aHP sp�otplugN�S�p��O�-inb�S/PPG ��0~�r�C(SC�P`��LC���J�\sw'�� � �� t����^ |���trsv\���1.pc
���  fx_�2����b%3��B	4.:�B��5���&6�#�C7�	��B	18���Btn
�0���=�F�n��sN�N�omi�p Posei�Q���NN䀇549~�Ї�`(pB�ѝ���TXP5
�n��os\nmt�p "NMTX"� #1�П]�e9t6�OMP�.�����-fxuif�N�-fle��b�F�XUFd�Ё�*"(�'�6	"$  f !"*!�sq&_�е�o$�	 ,]�t#w斠rl�o(uf.�vr.��'
@{in�cus.��3&#2+1��"��M?U4 K?]?�?�?�?�?�?�? �?�?�?O#OPOGOYO �O}O�O�O�O�O�O�O �O__L_C_U_�_y_ �_�_�_�_�_�_�_o oHo?oQo~ouo�o�o �o�o�o�o�oD ;Mzq���t����� ��	 {  7j$���v�|��r�q�j8�47\wti�v ��/���a��/�q���weW ��=���{47,r768R��asyArm&�f�un?�f�C�R� �S01h��Ь�(X�t E����X'��~�\popupcAt�#Ã,��aN��M�-Shelld�R533R��J�/ (Mu��-[����;'���vrdb�c2
5C�%� �enoio.fC�EnH�ced I/Od�"�3���J�6v�ŗ�p��ܷ���repa��c���?�accu�airR�AP�AirS�6;�0�kz� (\�p���O���S��ca
���4�O� �2��!S�� 2 Gu�c�����49 R63z����(������@��g�aΠib�#A�oSEL�^�/����!C�`�n,a�flowL�3� AF-AS-FMS��mmP�AFSM��x�2~勁����(�غ����S�˴��afgl
2��G˾!��P̴ۢF�̳2V�F�e�AFް��������᳣�O/�e�2�ȡ̱��d�̱2NL�AF2�Ͻ�2�� ���l��RӋ1B�@sŚ���x���!w��P��G�_�ɶ3��A�!㹽�AS ��~�5� �����`#����v�LO��.���˱������C�clrpt�hR�ic Cl�[���thϜ778ʪ�7��gv�ȀBas��@����� �ᛲ���>�S��㒐��tpqe=���s�sub������n��=�� /�w�set�����"�q���w�q�Off-�line Svu�lari6�>�85x>���[�85 ( ���tya���sia�d\tp� "SIAD�/���x�,k�plug���Dispense� P� j�=�SPL%G. 9s�(����g-i��� ���e�a�\sldsp�i�"�U8���0� }L% Trk F�� ̀<��>��ꖇ%\���For��tq𻠏(�]tcyc� "T�����k�tGgtp�/��!l��la��-#ptkmisc5#�"!�����w� ~��os�able EOAT<�_�G�����(@��
� ��3Q!b��"t���%1��Fou���os1�)t�47y
���47 (U4��on�)0�_�K1�2�+3��7��a�J5��r�70��ervo �Tip Dres��08>���0�ȁH7�r7��A\turnd @b���`D�'�����MHb<+�2	��@_��Lq�32]?C5/�S��A�in`�� ���'gcYht ��VG��r��SGCH J*!J�643>�Q��GN� CfQ��cT\s�vsvch��CH�/���TglgouV/�[gnc]���_��P�R�	dV;�sgd�ia�Ssb co�rey2XDG�P7!0�P�Q{<�b(~d7�p`O��rc�cinib��^btdw�j952�Ҵut@unSC9S<���R Jp�iH8r({��u����q�Pat݂c�w������ux�h8�69I�7�l�

/F,
1v���3� mtsv "�MTSV�X�j983\R���&P��s�ov��&_p���vruk%_c6�� 8����pex_�r�col$Q����v��v"�r���&�sxcM.Tool��k���=MTOF7p8�4 J571 R�814�!7E�ǈ�(��q���	mtofs�0��ߘ�2����pt�a��lle�to���k�PTLC��9����J9�813���H���T�4��9��`k{;��1�a\p�mk920 "K ���S!R����1�Ȥ<���2¢2�_�ި�4���!�ڣ�a6�1¡4��0����E�(ܣ�q8�4f�4C�c&0�5f�����ݤ��9��7f�7C��ަgr~@"GRIP".��쿶��1i "OP�TIC��1ݧpalf "PALF�Q���@�{ĻPSSU�C�F!ަcpt "U�NIT�S7mަxf�XFER��ԃ��et��L�U�&ʾ|ŏ��psysdjଭ/����mޤopti��Kޥ����7߹�ssu��+�ޤcpG!�W���er��S�N�t��ߞ�sӸ��d+�[�a�dpՂzaAdap?t CtrlF�3q50E�G0汫�_|���l\apa��R.�C����a�1l"�wgui� GUI��T���c[�c��xogJoU eWtra�&��u��f�86F�� (��b�r6��re���3�ETN;���S��X��5x��j7�22\cust_�wv6�RS�v7x�RS�[8�;QU	�9�KUwv10|2oRwvpat-x�T�ange/;xUh`#C j80��WeldCond#Mo���H�JK�#7a�Dq (T���i~J\atk30e�`��R�1�{�wm]gMON�_�0\�@$�_��$Xg��p� �b��"At��%stop�/rù����Zd��y8N4C�ir��ld Pr��XvF�ׁ��K���1��cS7�O1�1�\q�-\?8�at_ufrm.� #ER��7xcArc Ab�nr�l \ito�b9  �H552}�121� [prc��2� a�1AAV�M ��20 ���J614��@T�UP mch "n#@545�PC#B�6��VCAM� awam�0CRsIMe_@UIF��n#A28 0`vr_@�NRE�b.@R63�1�s�0SCH���DOCV li{si
@DCSUE��#A045pR51EIOCe t��0�542}�R�A96� pC
@ESET5 ��c
@J5K@���#@7K@;bMASK acryv@?PRXY cw1wBy7%��0OCO P�ht�B3�s;B2 � Q�B0�p pa�#A@4�;A39�0F�o�@H^SI�L�CHK�@59�@O�PLG ��;A03y ��PHCR :�~PCSP  GW�f�R6 ��;A54��nPDSW@_f�0{MD;P "FO�@�OP;P�PPRO�!ÏB7 mfor�k�B0�UPCMFt	e�@4f507�U��@5-hg��!fRS�T-f69`clm�PFRD@�SRM{CN	eH930�e�SNBA�USHL�B	eSM�`mex�te�B6�fPVC�-g2�`��~QTCP��UTMIL	f78�95@ups�`PA�C�fPTX	eTE�LNrd�R9Ef8�@w1 mpus�h#@958Ef95�7	eUECKYuU{FR�fVCCM	e�VCOR	�k.v�S@IPLU�@I ���_f�qXC k�Z�_@VVF �?WEBP Y��a�TP��t.�pR626 T Inp�CG�pnF�I�=� ��6�PGS��R3_q95 71�8 P�0738 �f��1�@
  ���AC`6�A63 7�94�B523�5R�65�1Sua553 ��A4�@gC=@�1qED064 tamapF���O�6 sths._@/LIO ��w^p���5 - HefPC�MSC��ӂP��5}1@STYL t��_@TOP ��PR}5{@Wave,�P�RSR ��A80�1UOL�Ph� v@O�PISY0��`� �w.��0L�p}��St��t^pETS��fun�0SLMT�Y0��B9 623��A�`E�5FVRCx�0_��NL tj�Nwp001E��2Er��3)E��6 j��F:@U0'@BDݐ5ME�ݐ8 a֐��U0@�`6������5�󔫑?@s@S���0Ff�61�=�3 ��l;��@69�U5`d*�faF�_�7 ��݁a�8Y�04^�9���_�_PT�up��2�0w0��6u���7 ����@��8 �"��9Vu�us�0U�1aw��㢸�{@Ʀ�@Ҧ33bݧ38`���`
�@~�7 R.$M��&/�K ���9����40E[�1̀SeԂ@]�2��Ea�AN�RSل� �334A���拰��n�e���Roboz���ne�t�����ደ�9����!拰j��\srvo���4�@h��p��x�����Srv��_t ROB:PM'��e�4��5��G�n�rr��b*ŋ�ite��ӿ�5�-���6��s35v��564���7@Main��tatio����6�� ��������o�ŋ�S��, '��� 溋�\��\cc�� "TORC���������L��crV�C�R�����5'�xk965������N���MО�6�����;���o_��w5���0�ch��y6���v.j�k��iw2��
���x5�����2. ���n���3V�h��z��5���uif����c��_�3E@H���,�l�����T�1���T�2�(�Z�l�4z���?������/�l_i��}3Ѧ勰�0� |�=��  Y2?��jog\djui����og��awm�fr� f��F� i�us�� Eq LibJ��6K񄐞S��/3�� (�b, ��2�7�_5'�\���� "MF�����
d5a��n7y57eM��mK��߽Ҡm���g ������̞At�w1������tw����#���6 ink��0LR .��6·�J852���J5�97�98��88�J�!�1^%N6��b��GN ��k\etl�@.�CO���O#A>` "ALNK
�>�%rd_�PB�� �"\wr*1O=�"�lS ��P$d��08�8����PN ARC��PRM�3��B� �0��Nŋ��!8^����1SU P��$P��Ç�H���0��p�>�3mpana/'��8�0�1��H57X��85n�����ã0 K�BH@��<��1�Gbel������R��<D41��HDY�dhen��8<A��ȄD���Cm���EN ������D.��E�ن!� kemp��D�4�3�m:re�2�r�pEf"sFMIG�A00��37JR��P�>!�IGC (�P.��E�%�чߑT� av�s��IGE��G�m�igco`'�mn�&NA�ц�favwavtj�VTPo~/lfrm "S�plGoYmsy�ASYqo�/lpdhV�PDH��oYktpdl7�D�L�o/lrf�`CRF�d�y�p8�3b���s�`.vr3hy�rLO5ccr��p� 4c�§��q��� ���������R�R�S!g�S����.�o��.�x�Z=fArbt\�`�c.2  ��; _	b��! TertiB�
ELS�P�2�Ug���YL (Com�myle seDU�%)��bգ�s���'�ps01 "P�S��.#le\pscol���u.т�ry�Pr: ��v�ׁ�Q�4syrsr���-���ice �Requ��g%��S�RS�2K�9�P6455.�9R S�"|�$���(����vb��/h�,M�ۂfO� "��s�O��sr����D�aP5A��+�m����2813�P�49Z�89���A��{��Z�.���g�st�M�\����|�
?�M�utl�v�'��&Q�N����q sp�dramj�!�pe�ed.�pf%�Q��NsN05���J67�2�NĻ�� j�(��d �RH�-�	D��b "RMTX"��ƏE��  ;�2 "S�0q�QD����slmt�of�t� mi��SL���H6Q64�H�62F�20�60�7B��P�38e�2C Hk�e�s�;�5l��62K�79��79�5�79��609�j�1F�1x�4��5���2����H6��8�43[�2s�825j��6�MT+�"�봠�6����f� �"����S��\f�봆봖�0n�-� Positio�l��esf 봷1#N1h�ݻP(���ti��,봥�ǀ�v�n1Z�POSs�� �0� �h8�73�r�rive� Axes+�H8���4di��(Du_al Dr�sΕ$�Ȅp��C�\B�j�`.�kŔ*�ex�s�j� De)�1�6�3����AM Indexjź��<�&�\ami:�ṡ �mi&�8�ca��sC��nt An7gle+�CO;�����봗#COM��Mom���������ggou���! ���
fl���Env�i� m���6k�d�8c20)����fl(�<2� |�r�봇ionΓ{�ǅK�r?772\ic��$(	� �x0Z˱;�:�2atzn������c�TJ�yncIsns�p��R76��� �#���Xj�rm�SB����T�b5mK�masyA`jբ�nc\��MAS�Ir�{��ba�s��ulti-A�`�6V��7v!� +Ռ�5k�NN�P ��s�e��!\��FR�LK��v�k�h�dzՎF봅"frlIk��&�m
ŊTr���C��il/-&e��r7��0Zon�d ��:���� "ICRZp�%Qg8��Piabic..T�IAB0c���0o�e�I�0V�E �0��1 (�1�4��0`濡�0�C�2\i�0t� IA˱����"\�@AiciAC�0�b��!�1�1��!�0m�ain�sDP�1n� C7`[��0e�DL�PV�2�0��hpV��P M_@��̘��O]B�ưI:A��Єdp�CD�O�F
"�0N>I�A�B��H�0_�Fd%4�eo@nn Stan�A|[�'"� MCN�6>�90�096:�s�A5j��0�Q=���H�0����Q�2~Q(Remx^PkAeSdardI0࠸W2�NQ�0\tp�rcmuǰCMU��ku�1�TRP\rc��0�q��jBRSUF1783 �0uip��[�܋Ae�J61S 59�Q�I�0taV"i Eq[A��Ζ�Rǅ�!ȡ�jt`�Pcp��E`sr��A�Qvb2 �Q4⦷ka�@xa�0#��-���1 �a:��1 awmgenl�qޛ0ener��We7ld zQiboX�0�AWMG�U7{o �_q(G>t�A�`%�b �;�d�60t[A3rt�1x.y�R mshcq@|�3��n she�qxqGR��1CMSC�U �A���RhjQ����p��0l�0rd$�1�8 �p[a��u\qsh�� PSH��� X  ������0   (L� r wKq�1/F�e$�Q7�Ij��\cl
A "J����0v H\j�Qcle��C"E�S�Heӄuyb�U��`{A�ybmd�prm"�8�zali_varsS�����iconu���db�g"��0Iz�ցrgpged"��1�&��� Ԅm_�0�1�i<�Q҃m102؟��e_no��ȕwr�spq����wrp�irS�[q>��0ga!s��Y��1��_s���cwr������ffӯE�inch30U���extwd���'wrc����'�DՂrdS�Q��0!�i�����aN�b�i ����0�Ə(�/i���RF�p
q���saj�c�a��ntKCMAP	 ���O D�B�)�T��f�ap"Qj�APCp��Z���0stm(P�STM.Q{� ��a?pcevre*a�o��in
Au7a*a��is
�rbCISD{ G�QMete/`�3�0T56��i<�pcQ��Q7�ar >��,KQ�Y��(�\sl
(�gr0S�14�e���q�	B..i�A�����d��/�[a��>ֻ1��PQ�d+Q�G 
�(5���M�Q�O K�џ�` +�2�`KQ�����B��Kq��GT��sU�0ӛ0�S30le Act��C�8R��Y
AQ�4�.��1�㵏�I��\J�ds��SU^�%����{A�#���s�!j�691.f�1Se�rvoTorch�9��6Jv�K� 91� (�K�A���Qs�vt��VR��AR9C
�es4 F���Q4��MU�dq�v�z�vt/���5�+Qt FEv� ՛0"S`�0�h for Alwumi��982��� 82������ ��	��d�{���oo�q��l��L��ϊ��\srvt.vK�3e��0�hP�AS`�� A��<
�/S016F�85��0�*�(!ez���hS�ATNQ���h
�0"P�QNG��	t��2w�ADW����t��ҋ����wenmr�8snh�anced Mi�r�bmag ��bR�69�Q90�+�E.'KQ I>!��I""�\mjQr�MIR�c;� � e$!.b�0�6b"%�tmbust�cpy�Mod�  TCP��REˑX �nvkAd�8���!KC�P>� \�$�Pm>:1"MBUI2���i2d0� i�+�%��p��930�sPROF/INET��OJ����J93+� �0 (��5��>鋁Y�3�Ppnio ":���xp�1"P�q(@RIO�/�ǖ$A��u�3)tj96Od:��@gT�UHc�67J�O��Q�`F�SW䑡@���?K67\fswpr��qW+F�}�A\f_�a�ch޷	�A;ber�4���96�p_fw�d!6���f_re�a/T[O 'Qneu4��_�Rr��sR��C��Qurn���%Seinא� $Ssw��t�_fswcol��#�n�AQ��Ak�c�vvcuj�2�iRCalib Vz!�nc Utl4�V'CUT� ��1?�b�(�a��VisFu�cj���`k�vcc�U���c�tpfi a�_z��`p6b�_+�apset�3���c\z_�p{���k��u�KA4���c��j98�8/�To��ors�1�!�p.�=8�? �p ^ol +!�8�+��p\gf*���D�sT�c���VM�as@��9�;� |ë����1� Po�sij�����ord`t���v�
�02\���up޶�����r_Gdc1$AB�As.��I[\N�bjA n�e��b���򾿮��ۿ]���+�ޘ�� _ywQW�� k_c0!y�t{G���F4�1�k�nifi3 sp)eY��94� a�1�UI n���v�>�k1|��`�\frco���
�j9��1�Br�ake ch:�fP�`0�{Q�5GJ��(�ck�rpȺ���˕51��b��BRCHUCD ����P�����5/�C����mulaneous�=l���>55`�loH��SiɀST�D u�LAN�G ��!�cs���0C�T��\c�scsm���1 ﳔsﳠ�=��C���N�dss' ﳣ@gc S�F�
�`����3�V68�ςF�,��sﳥ�s\��u�ߣ�ć�N��r69����gno[st�eo� n�@����1�U�i-� �9��C�ﳵ�7�!�=\�"DVMV�����"r6�Đ��!A !��p��U��� tr�D!ﳆ�Q2ﳡ�[�4� Tc�����er�!��q+�\pc3j����܈Ƴ075.�os.Re���rN���g� �2c�6��ė�� ��Ͼ��75\pt�TJC6���b������@�Bg�ė@I>�eS�i>��80�oJ979a�08 1X���(Iepi{�UL+�oﳔ#�a�~�f "NRU��|¡�prsta2�|£��gutl.���RBT��OPTN�q0\?�r?V�@H nr?�rovq�?l rb?r�DPN���!�rrGdfi���u�����basic�ߡ�fc� �J�Ġ�A-�q��H8C29V �$��9�@@������Ph�c "F2�
Ӡs29���j83��ެce C�to{ur� UPDT3³5����Fo��on���a��Ӵ�Q8�hof�f���r� 35�fnV���r���\f�V�����\fcn��rg%3(��% ��r�A���@���6�%�D� E������g0=� �$���$n��/J1!46%u��C/ T0�\> ])A��av2t�p�0ޖ�0v�0�2v 6`�0���0?U8�0�1�Br�0���0�4U0L�vpofs`1|��1�3>y0� mgp�s�0Nv�<un�Q�,x�0�4se�5ҌBT0��b? cellf�1��el�0Cp���1���R�1�f�B��519�1ll F�B�0��p�0b�C�Bn�0fncl��"RA��Zx�0^V�Bfndru�<�AsIND"�1�>\�A�1\fn��t�A�^f�0t�B&PTPex@jA�?�@�0%QTPc�1�v�1u�B&Ptqd�~_�[ Q�2�V�Gj�7��0- V-5�00i/�010i 3D�0�[S���15�`ab`�13�DE��0N��<9\cGalc@�_.27�0?vsfit3Ep�0�{a���07�u�0`.�`Tra�0B��K	J�a�MJ�`�b�e�1��bE��10Ov�0j�`\que�1�?�3FArpo��8_�`8�1�epush3�� H���0}s\�М�v��/�qkm�1ޕ\�s�wa�?�h�qain<j|wkclb*O���?qvs
AJ\uds�blt���een�n�g�|wigchik��uv�avuA��s�� |�{�0  �0тv��3��_p��FA���GA"73�1cr�o����,�v�Apo ��0�8�a�jB���iR�qon ErSro9���.m�FQ�A757�Aж�1��� (iR�A���R.�]kZ�<d\mherhd�AH4P���}��\ire:AR���ree���/0�B@����l��Z�h:Ahd���� ������j��c�v�a���`�1SP �APAS�A��SAS�z�09 �q CTsAMڠQTABڡ5P�AGz�13�Ҷ�Π(�`�Q����px&u/M��pas\�aama�s+�=�
AF�0�c��s��bia�B?�����VS����VSIAС��D�q��Ⳳ(�A��vAC��  �6� �����1 � !   ���� �Ó0(�8 ��\���ұ�(H� ��]ia\ia�`�a�`�4��P�g�QoiZĳ|�c������ � ����*SYS�T�EM�0A �����$ˢ��S  ��0����������ATSTKSIZ�������0������ +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy �������	 -?Qcu��������*������TART_T� SAG��$D���IGNAL���SARTUP_CNfQ/a/s/�/�/�/��/�/�(J�2!
�
 �/??)? ;?M?_?q?�?�?�?�?��:99�$K���$FEAT_�DEMO C�����1@   �8MO O MODOVO�OzO�O�O�O �O�O�O_
__I_@_ R__v_�_�_�_�_�_ �_oooEo<oNo{o ro�o�o�o�o�o�o A8Jwn� �������� =�4�F�s�j�|����� ��̏֏����9�0� B�o�f�x�������ȟ ҟ�����5�,�>�k� b�t�������įί�� ��1�(�:�g�^�p� ��������ʿ��� � -�$�6�c�Z�lϙϐ� �ϼ���������)� � 2�_�V�hߕߌߞ߸� ��������%��.�[� R�d�������� ����!��*�W�N�`� ���������������� &SJ\�� ������ "OFX�|�� ����///K/ B/T/�/x/�/�/�/�/ �/�/???G?>?P? }?t?�?�?�?�?�?�? OOOCO:OLOyOpO �O�O�O�O�O�O	_ _ _?_6_H_u_l_~_�_ �_�_�_�_o�_o;o 2oDoqohozo�o�o�o �o�o�o
7.@ mdv����� ���3�*�<�i�`� r�����Ï��̏���� �/�&�8�e�\�n��� ������ȟ�����+� "�4�a�X�j������� ��į����'��0� ]�T�f����������� ����#��,�Y�P� b�|φϳϪϼ����� ����(�U�L�^�x� �߯ߦ߸�������� �$�Q�H�Z�t�~�� ����������� � M�D�V�p�z������� ������
I@ Rlv����� �E<Nh r������/ //A/8/J/d/n/�/ �/�/�/�/�/?�/? =?4?F?`?j?�?�?�? �?�?�?O�?O9O0O BO\OfO�O�O�O�O�O �O�O�O_5_,_>_X_ b_�_�_�_�_�_�_�_ �_o1o(o:oTo^o�o �o�o�o�o�o�o�o  -$6PZ�~� ������)� � 2�L�V���z������� ����%��.�H� R��v���������� ���!��*�D�N�{� r����������ޯ� ��&�@�J�w�n��� �������ڿ��� "�<�F�s�j�|ϩϠ� �����������8� B�o�f�xߥߜ߮��� �������4�>�k� b�t���������� ���0�:�g�^�p� ������������	  ,6cZl�� �����( 2_Vh���� ��/�
/$/./[/ R/d/�/�/�/�/�/�/ �/�/? ?*?W?N?`? �?�?�?�?�?�?�?�? OO&OSOJO\O�O�O �O�O�O�O�O�O�O_ "_O_F_X_�_|_�_�_ �_�_�_�_�_ooKo BoTo�oxo�o�o�o�o �o�o�oG>P }t������ ���C�:�L�y�p� ���������܏�� �?�6�H�u�l�~��� �����؟���;� 2�D�q�h�z������� ݯԯ� �
�7�.�@� m�d�v�������ٿп>��  �� $�6�H�Z�l�~ϐϢ� ����������� �2� D�V�h�zߌߞ߰��� ������
��.�@�R� d�v��������� ����*�<�N�`�r� �������������� &8J\n�� ������" 4FXj|��� ����//0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O �O�O�O�O�O�O __ $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�?��?�?�?�9  �8�1O(O:OLO^O pO�O�O�O�O�O�O�O  __$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv���� �����*�<�N� `�r���������̏ޏ ����&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ���*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�?�?A@�8O,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o  2DVhz� ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟ ޟ���&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ���� �0�B�T�f�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p������ � ��$�6�H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я�����*�<� N�`�r���������̿�޿���$FEA�T_DEMOIN�  Ā2������INDEX�'�6���ILE�COMP Dw���h�5���^�SETUP2� Eh�r���  N ��[�_�AP2BCK 1�Fh�  �)������%����� k���/����[���� ߌߵ�D���h���� ��3���W�i��ߍ�� ����R���v����� A���e������*��� N���������=O ��s�&��\ ��'�K�o ��4��j� �#/�0/Y/�}// �/�/B/�/f/�/?�/ 1?�/U?g?�/�??�? >?�?�?t?	O�?-O?O �?cO�?�O�O(O�OLO �O�O�O_�O;_�OH_ q_ _�_$_�_�_Z_�_ ~_o%o�_Io�_moo o�o2o�oVo�o�owɺ��P�� 2���*.VRN�`*Qw�c}��e8p�PC���`FR6:��~�"��{TF�F�X��uC���)�x����f*.F;Dُ�a	�sǏ���<*���STM J�S��^��pK����`i�Pendant �Panel����H ���p�ϟ���3���GIF=�g�r�S��8"�����JPG����r�ׯ����;��zJS�E�n��`�\��%�
JavaScrgipt��ůCS����q�߿�� %C�ascading� Style S�heetsϐ`
�ARGNAME.SDTMϰlu�\a��ρ��Ģ�N�	PA�NEL1����%@u���%ߜ�����2߀���n�+�=�����3 �����߯���V���4"���v�3�E����Y�TPEINS.gXML��}�:\�������Custom� Toolbar�6��hPASSW�ORD��nFR�S:\y�8� %�Password Config�� �o����9�o]�� ��"�F��| �5��k�� ��T�x// �C/�g/y//�/,/ �/P/b/�/�/?�/? Q?�/u??�?�?:?�? ^?�?O�?)O�?MO�? �?�OO�O6O�O�OlO _�O%_7_�O[_�O_ �_ _�_D_�_h_z_o �_3o�_,oio�_�oo �o�oRo�ovo�o A�oe�o�*� N�����=�O� �s������8�͏\� 񏀏��'���K�ڏD� �����4�ɟ۟j��� ��#�5�ğY��}�� ���B�ׯf�Я��� 1���U�g�������� ��P��t�	Ϙ���?� οc��\ϙ�(Ͻ�L� ���ς�ߦ�;�M��� q� ߕ�$�6���Z��� ~���%��I���m�� ��2�����h���� !�����W���{�
�t� ��@���d�����/ ��Se����<�N���$FIL�E_DGBCK �1F��� ��� ( ��)
SUMMA�RY.DG���MD:!a� �Diag Sum�marybo

C?ONSLOGW:�L��tCon�sole log��n	TPACC�N�@/%(/e/p�TP Accou�ntin/o
F�R6:IPKDM�P.ZIP�/�
�/�/q� Exception�/�+M�MEMCHECK�[/�Pq?�Me�mory Dat�ar?ra,])>]1HADOWg?L?�^?�?�3Shad�ow Chang�es�?�-��)	FTP�MO�?�QO|7�mmen�t TBDzOr�=t)ETHERNEToO�01�O��OtEther�net �fig�ura?udADCSVRFnOTOfO_�1%DP ve�rify all��_�10"�?UDIFFw_]_o_o�0�%�Xdiff�o�W01DPCHGD�1�_�_�_�o Xo�o�S!�Gi2o8foxo �o4�oGD3�o�o�� #�GvUPDATES.�p���FRS:\���uUpda�tes List���PSRBWLOD.CME����Y���PS_ROBOWEL�Omޏ �����8�J�ُn� ����!���ȟW��{� ��"���F�՟j�|�� ��/�į֯e������ ���T��x������ =�ҿa���ϗ�,ϻ� P�b���Ϫ�9ϣ� ��o�ߓ��:���^� �ςߔ�#߸�G����� }���6���/�l��� ������U���y��  ���D���h�z�	��� -���Q��������� -R��v��; �_��*�N �G��7�� m/�&/8/�\/� �/�/!/�/E/�/i/�/ ?�/4?�/E?j?�/�? ?�?�?S?�?w?OO �?BO�?fO�?_O�O+O �OOO�O�O�O_�O>_�P_�Ot__�_�_  �$FILE_�{PR����P����X�MDONLY 1�F�U�P 
 �;_o__6o�_Colo 5_�oo�o�oUo�oyo  �oD�ohz	 �-�Q���� �@�R��v������ ;�Џ_�����*��� N�ݏ[������7�̟ ޟm����&�8�ǟ\� 럀���!���E�گi�����ZVISBC�K�X�Q�S*.V�D�a�ϠFR:�\0�ION\DA�TA\L��Ϡ�Vision V?D file���� տ������/Ͼ�@� e�����ϭϿ�N��� r�ߖϨ�=���a�s� .ߗ�&߻�J����߀� ��9�K���o��ߓ� "�4���X������#� ��G���X�}����0� ����f����������U�ZMR2_GR�P 1G�[��C4  B�> 	� �Q��� E�� E�@����`
� OHcGP��K���Jk��?� `ޙ :G:�<9{�H�A�  �dvBH�C��=N�B�ƈ�`��� z  D����>��	@UUU�UU�`/����#@=ud�ѽ��H=���=�~�=�y�C,���;��.;!�9����:�b:�l�?��/ /�/�/�E�  F,D �!D�`�#�u�-���E�� �!D+��2C�dR_CF�G H�[T ��/O?a?s?�NO� �X�
�F0�1 �0 � � �0��PRM_�CHKTYP  ��P�> �P�P�P���1OM�0_MIN��0<���0�P]X�PSSB%3I�U�P�#O:�CCOUO�UTP_D�EF_OW�P:|�YpAIRCOM�0�{O�$GENOV_RD_DO�6�Rn�LTHR�6 d�E�d�D_ENB�O ��@RAVCxJGC� ��[OF_�/j_�x_�_7�P[�QOU{ P���B�8�(�_�_�_oo/  C�f`\Vo�X4�oYm%~oBȽ�bp�	�Y\OPSMTS�QY� @ed�$HoOSTC%21R9���G�  M�:}k;8�  27.0�p1t  ek�� ���z��1�C�U��x|�	�	anonymous|�����@Ώ��7:� ���� ik�P��t������� ��������9�ӟ ��^�p���������� �+�-��a�6�H�Z� l�~�͟����ƿؿ� �K��2�D�V�hϷ� ɯۯ����#���
� �.�@ߏ�d�v߈ߚ� ����������*� yϋϝϯϱ�{��Ϻ� �������Q�&�8�J� \�n������߶����� ��;�M�_�q�F���� |������� 0S����x� ����K!3/G i/P/b/t/�/��/ �/�/�/�//Se:? L?^?p?�?����? 	?�?=/O$O6OHO�/ lO~O�O�O�O�?YO'?��O_ _2_D_�bqE�NT 1S�[ cP!�O�_�R w_ �_�_�_�_�_�_ o�_ ,ooUozo=o�oao�o �o�o�o
�o�o@ d'�K�o�� ���*��N��G� ��s���k�̏������ ��׏%�J��n�1��� U���y�ڟ�����ӟ�4���X��QUICC0e�A�S���w�A1�������w�2����T�!ROU�TERU�1�C���!?PCJOG�����!192.168.0.10~�~s�CAMPRT��ѿ!�1��ƃRTn� �2ϓ�YTN�AME !fZ!�ROBOϛ�S_CFG 1RfY� �A�uto-star�ted�4FTP�?,��?�OW��?{� �ߟ߱���hO����� �@�.���e�w��� ��6��)���=�_� �F�X�j�|�K���� ���������0B Tfx�?�?�?��� �3�,>b t����O�� //(/:/����/ ��/��/�/�/ ?� �/6?H?Z?l?�/�?#? �?�?�?�?�?K/]/o/ O�?hO�/�O�O�O�O �O�?�O
__._QOR_ �Ov_�_�_�_�_OO 1OCOE_*oyONo`oro �o�oe_�o�o�o�oo �o�o8J\n��_ �_�_o�;o�"� 4�F�X�'|������� ď�i�����0�B� ����ɏ���ҟ ������>�P�b� t�����+���ί������T_ERR �T���"�PDU�SIZ  ��^�ɐ�9�>R�WR�D ?�Ō�� � guest��������ȿڿ�쿣�SCD_GR�OUP 2U�� U����1��!���2�ǒ  ,C�	�$SVMTR_I�D 2�Ti��$GRP_2�$A�XIS_NUM cY�z�f�NF���SV_PARAM�iɑ� ,$M�OT_S��TTP�_AUTH 1V�1� <!iPendan���J������!KAR�EL:*����KC3�C�U�+�V�ISION SE!T��ߊ���!�߸� ��(������e�<��N��r����CTR/L W1��谡�
��FFF9�E3�FRS�:DEFAULT��FANUC� Web Server�
��z��� ������������� ��WR_CONFI�G X!��m��"�IDL_�CPU_PC0�氡BȊ�K  BH�1MIN<)�OGNh�O+�`���7�3 �NP��IM_DO���TPMOD�NTOL� �_�PRTY�K�O�LNK 1Y1� ��#5GYk}��MASTE� ����	OSLAVE� Z1����O_gCFG��UO��|��CYCLE���*�_ASG 19[l�
 ]/ o/�/�/�/�/�/�/�/ �/?#?5?G?�0"���`�5�_��IPC�H/���RTRY�_CN0���SC?RN_UPD_���9� ���\�1�&�O&��$J2�3_DSP_EN�B�01�%�@OBP�ROC%C��JO�G�1]1�8���d8�?��R;�OR??U�S��LQ �O�O_#_�OG_Y_k_�}_��'ҟ_[CPO�SREEO�KANJI_�K��S1��3^���U�_�UCL_L[ m2�?�P�EYLOGGIN��&��}A9���$LANGUAGgE m��*� �a"�LG�2����V������x&а�Pi���Q ���'0�������MC:�\RSCH\00�\�}`N_DISP `1������O��O �LOC�BD�zj�A�cOGB?OOK a;+~@°���q�q�pX Cy�����*�=�10�O���	�u�y���Fu����!ua@BU�FF 1b ��2��ڏ�r������ �$�Q�H�Z���~��� ����Ɵ����� ��M�D�V�����DCS� d�} =���L�����!�����|!���IO 1e;+G 
OZ����Z� j�|�������Ŀֿ� ����2�B�T�f�z� �ϜϮ���������
��5�Ez TM  2{d�_c�u߇ߙ߫� ����������)�;� M�_�q�������qw8�SEV�02}.4�TYP@�R�3�0E�W���QRS? Ko|���2FL 1fC��0�˯������0%7h�TP_`@��"�k}NGNA�M%D�e���UPSF*pGI�5a�5��_LOADB@G [%2z%�1D�U>MAXUALR�Mm7�{8�_P�R�4�0�sM�C-pg;)[�q�s��Pc@P 2hVk ��	"���0���t���� � /ɨ/O/:/s/V/ h/�/�/�/�/�/?�/ '??K?.?@?�?l?�? �?�?�?�?�?�?#OO OYODO}OhO�O�O�O �O�O�O�O�O1__U_ @_y_�_n_�_�_�_�_ �_	o�_-ooQocoFo �oro�o�o�o�o�o �o);_J�f x��������7�"�[�D_LDXDISA� B�3�MEMO_AP� �E ?��
 �c���ɏۏ�����#�5�ISC ;1i�� �M��� �b����L�՟�����J�C_MSTR �j���SCD 1k����g�韋� v�����ӯ��Я	��� -��Q�<�u�`����� ��Ͽ���޿��;� &�8�q�\ϕπϹϤ� ���������7�"�[� F��jߣߎߠ����� ����!��E�0�U�{� f����������� ���A�,�e�P���t� ������������+�O:s	�MKCFG l'�n��LTARM_�m
���q��|�,METPU9�d��/�ND�CMNTd�% � n'�c��{|�%POSCF1=<PRPM0�STOL 1o'�� 4@C�<#�
�n�/'�/ /1/s/U/g/�/�/�/ �/�/�/?�/	?K?-?�??�?k1%SING_CHK  �^t�ODAQ�p��=���5DEV }	'�	MC:�<�HSIZE��C����5TASK %�'�%$123456789 \OnE�7TRIG 1q`��%H��OA��O�O�O�)�>FYP)A�E�4��3EM_INF �1r� �`)AT&F�V0E0�Og])�OQE0V1&A3�&B1&D2&S0&C1S0=V])ATZg_�_�T�H�_�_vQ�Oo�XA�o?o�_coJo�o�o  M_�oq_�_�_�_�_ <so`r%o�Q� ����o�o&��o�o �on�y3���ȏ�� �����"�	�F�X�� |�/�A�S�e�֟���� 1��0��T��x��� q���a�s�䯗����� ,�>��b�����A�K� ��w��ǿ��ɯ:� ����#���G����� ��ϡ����#�H�/�|l��?NITORL�G ?K   	EXEC1j���2��3��4��5���@��7��8��9j��6������ �����������Ҁ��������2�!�2-�29�2E�2�Q�2]�2i�2u�2���2��3!�3-�3��һ1R_GRP_�SV 1s<[ �(s1@ʾ�L=��-k��׮]�S��=FA_�D�,N�PL_N�AME !S����!Defa�ult Pers�onality �(from FD�) �RR23� �1t)4�x)4󭸬��0@ d p*<N`r ��������&8J\n�82 ��������
//./@/�2<�j/|/ �/�/�/�/�/�/�/?�?0?B?   ��\  � � ��`��  A_�  Bm0Tm0���0
Y0�]0�����  ��i0h0B�m0pm0�  C��0C�0P D��  D���2E@�2�2z�0�1�0 �1�2�0�9�2�0�6�4�EK  E+� E��6�2�0�2 A DJZ��3A@DI@�2�5�4�9�:�1;�7 �:�5�@�5�O�;�O�3ԧ1�1E�1��0�`� E���G�4E���C�@Q�A] Y$UP�5#V��DQL] hT�FQ8@�B UA U��T�R YU Q|UU� @�Y�Q�]�Q�Y�@B �YAP�1�R4oBg�U Xo�S�1Q`ong�Q�o �o�o�W�o�o�o �2DV`tU0DJ�xE�PE��R�q�S2O�  !l0��{q�d�sU0 ��}���tpI<Z*d����y����`q�0 b�[T� @�5?h0�p�T�?q�p�q�@uþ�5o���;��	l��	  ����p�XJ�����X � � ��, �ނO�K���K�zK��ɜK@0>KH?�K$�����О����5��N�?�{�P�@'�6\�����"��Iڿ��
��}v�����X�������0�
�=Âp¬0��� � >ڃ���#�^���l�Y"�0 ��q����͔��'���h������  �T��  ��`��v��	'�� � ��I�� �  ��-`�:�È��ß�=���إ$�@���Z����BZ��t'�5�o�N��j�  '��O��?��@�t˅@��@����X���B&d0Cf�0�pB�1��}q��C%
���e � W ��^�/�AB-`���$Ń�P� ��A�q��1ș_φ�o�p�πϹ� �
�`�����n� �x��ݱ�� ؀��:�m��q���?�f�f��0��� ���d�v�%��ߛ�?KY����|��(q���P�����ȃȄ2��?33�������;���;���;��D�;�$;�< Jl ��=�L�~�Z���=�?offf?��?&z�ޡ�A���@�,��j��u၄�� p���n���^約O�$� �H�3�l�W���{���`������+���F-� ��&��J��k��=,�ɘD�@����0�  F���� ��5 YDV �z�ƚG���/ a'/�N/�r/�/�/4�/G�A�0����O�tp��B�0h/?d/%? ?I?4?��-�A�0t2 -`|1�?�u�?\?�2;�<��Ŝ?���?�?hOO*�į��W*O�C��@�` Ca'O*�4��0�1�A���ܨ���C>�CR BA��Aˉ7࢙���"���z���q��=��\)xO� ʊ=��=qA�B)�{���O� ��(��g�/P�q�Bp���{���8R��K����J?&DK���	HwW�H�'���!��LA�L��9K��4HŀHH� h_�zP��Lm��J�sdHK� ?H-�A��_wO �_�_o�_%ooIo4o moXojo�o�o�o�o�o �o�oE0iT �x������ �/��S�>�w�b��� ����я�������� =�(�:�s�^������� ��ߟʟ�� �9�$� ]�H���l�������ۯ8Ư���G�$��� C���4�F@��8��u�8�V����������Ͽп�����?��F( Q�`���G� ���x�8E��Y��>x�	3Z�q_�Ϧϴª�����ϰ�fC3�g����̅��?�3�Ȭ�ـX�F�|�jߠߎ��5P��P������N�`����.���P�0b����7���
C@�C@5����
� @�.�d�������������������������&  ?JK  �@^���v�����2 wD�J�E����0��B}1q1}0C)�f@�AC@@�?F�C@J�m��C�����z���3��E�(��F���
/�/**@9$���4�C@C@���4�;
 */�/�/�/�/�/ �/�/??/?A?S?e?�w?�J�2��������$MSKCFMAP  D� �g!c!�>�3ONREwL  s��1��а2EXCFEN�B�7
�3�5AFN�CODJOGOV�LIM�7d@Bd��2KEY�7eE��2RUNULeE��2SFSPDTY���FE�3SIGN|�?DT1MOTWO�A�2_CE_G�RP 1zD�3\,�;_$�__q_� [_�_S_�_w_�_�_�_ o�_oPooto�o=o �oao�o�o�o�o�o :�o^pW�K�������1QZ_�EDIT�D�7�3T�COM_CFG 1{�=r&I�[�m�}
)�_ARC_B���DIUAP_C�PL��(DNOCH�ECK ?�; �������
� �.�@�R�d�v����������П����;NO_WAIT_L�Gl�	PNT1�|�;zi+F�_ERRQs2}�9�ф �����ï���3���^ńT_MOt�~{�x l\��D��8�?\_�I��b 6�m�PARAM:u��;�f&4����w� =� 3�45678901 '�9�K�"�j�|�Xψπ���Ϡ��������w��,�>�ѿb�ƃUM_RSPACE�?�R�o��ߥ��$OD�RDSP���F$HO�FFSET_CAqR�����DIS�����PEN_FIL�E��Ao����PT?ION_IOvO�A�;�M_PRG %��%$*t���WORK �W'C ���6���2���S���	� �a���6�C����RG_DSBL'  DCj,@����RIENTTO��0���2 ��UT_SIM_DC���2�2��V��LCT �P�����>��_PEXE���GRAT��\F$E��>��UP ���x E �/A'es	��$��2St)4��x)4����@ dRߺ�� �&8J\n ��������/"/a�2�R/d/v/ �/�/�/�/�/�/�/��<A/?0?B?T?f?x? �?�?�?�?�?�?�?������)P�  ��  �p�A� g B!@�B�Y�@H@�  ���@p�B!@p�!@�d�c���P �D�  D��NbBE@jB_Bzd� `A`@{A{Bx@�I{Bd@��F|DEK  E+� E��F�Bx@0kB�A�D�JZ�fC�A �D�I�B�ElD�I�JlA;eGJ�E<P�Ec_}KPs_aC[A{AEhA�m@?�` E���WxDE���S��@�Q�Q@�]�Y�U�P�E�V��T �Q md�V�Q�@�R�U �A�U@dcb�Y�U�Q0e�U˵@�ida�mda\i <P�B�i�A�P[A�b�o �g�e�chA�Q"w da4Bp�gx�� ����
����"�A @E�W���P�s� ��j�����(�(��� �O 1y(�Ho(�&��`�o0��C @�Eo�o��?|��C@�E��.�  ;��	lo�	�� ����p�X̰��q���X � � ��, �����H����H��H�P�uHV�2H�H_3��<���&��B�!@	�C����@�γ�4@L@�/
=�g��`@D��(�:�L�)�Aß�w½��ªV y�H@����p�ˣQ��֡�hD��D��  �  �������Q�6�%�	�'� � T��I� �  y��`R�=���x���(�@�������ʿ;��$�߯�r'�Np�"�  'F��:ą�Ca�B@CfBd�B�Au�G�Y� ��  ��C%�  ���^
��/V�B�`��p���;� ������wA ���^�'�M�8�qߨ��
�`��U�n� �x������ L����:O���Q��?�ffǏ���� z߶�%�ㅡ8��E�.S�?Y����4�|�	(����P���ő�������?333Q�����;��;����;�D�;��$;�< J!l�����6�޳8����?fff?��?y&2�A�D�@�,P�Q���-� 9�T�(���&����l� ����� ��$H 3l~i���� ��s������V���Dڹ@�U�@�  Fg�D��� ���/�/G/2/ k/�����-]/�/�/ =?y/*?<?N?`?��AL@��j��	�d�B8@ ?�??�?�?O�?B�'�A�*D�`4A ;O�0�?bO����S�}�?�؏O�O�O�O�Q��g��W�OC�>�P�` Ca�O�*�D��@�ALQ@I�	�b���C>�CR BA��Aˉ7��Q���"���z���q��=��\)0_�0ʊ=��=qA��B)�{�녨_�0��(��g��P�q�Bp���{���8R�MK����J?&DK���	HwW�H�'���1�MLA�L��9K��4HŀHH�  o�2`��Lm��J�sdHK� ?H-�A�Jo/_ �o�o�o�o�o�o�o %"[Fj� ������!�� E�0�i�T���x���Ï ���ҏ���/��?� e�P���t�����џ�� �����+��O�:�s� ^�������ͯ���ܯ � �9�$�]�H�Z���8~����KG�$��ſ� C�����@��8?�-��V��7�>�w�b���ψ�r������ϲV(xA�`����ϸ���0��ų�Y«N0߲S3Z�q_L�^�lҪ�x���߰�fC3�g��߶܅��?�3�Ȭ���ـ���4�"�X�F�EP��P��!�/���`�������`���0�S�>�V�7`�r�
{�{5��V����� ��������/I ��JXj�t��̪�����  ?JK  ���@.dR�r�2 wD��E���0�VB5A)A5@C)�P��A��@9O�X/"/2,C����2/�[/i*�CN�E�(�VF�i/�/�/�/R�*@�$�XxD�����O�|D�K
 �/E?W?i?{?�?�? �?�?�?�?�?OO/O�ZB��\������$PARAM�_MENU ?��� � DEFP�ULSE;K	W�AITTMOUTޓKRCV�O �SHELL_W�RK.$CUR_oSTYL�@�L�OPT��OPTB��O�BC�OR_DECSN�@{�N\H_Z_ l_�_�_�_�_�_�_�_��_%o o2oDomohAS�SREL_ID � +�x�@}dUSE�_PROG %�wJ%io�o}cCCR�@+�C�g_HO�ST !wJ!�d#�jT���o?s�qAs{�k_TI�ME�B�f�eh@GDEBUG�`wK}c�GINP_FLM1S�~�xTR��wWPGA � �|N���CH��xTYPEtL� hobo�� ����Ώ��	���(� Q�L�^�p��������� �ܟ� �)�$�6�H� q�l�~�������Ưد����� �I��uWO�RD ?	&�	�RS��PNeS��D��JOQ��TEbpF�TR�ACECTL 1���A ���% &e���� ߾��DT Q����ӰD ȿ 
 ��������Ď`!���
�	�
��0�B�hT�f�x�z��� � y�0y�0y�6�y��0y�0�ϻ��� ��C���C���:�L�^� p߂ߔߦ߸�������  ��$���;�-�_�q� �������������S�%��)�[�m����ã��£��£�� ��ң�ң�ң�&� ��£��£��£�~� ���£��£�£�� ���������	- ?Qcu���� ��������ߺ� �φϘϊ���� ���S_/q/�/�/ �/�/�/�/�/??%? 7?I?[?m??�?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O__/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}���[/���� ͏ߏ���'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߹��� ������%�7�I�[� m�������� ���!�3�E�W�i�{� �������������� /ASew�� �����+ =Oas���� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k? }?�?�?�?�?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	_Q��$PGTRACELEN  Q�  ���P�'V_UP �����VQ�^PBQWP'Q_C�FG �VU@SQWP��T9P�_��\kRDEFSP/D �v\Q9P��'PINnPTR�L �v]P8��U�QPE_CON�FIrP�VU��VQ�T�Y'PL�IDoS�v]�QEaG�RP 1�g����QC%  ��ᙚQA�=�qGY� GcX� Fg@ A� o D	��T	�P�d�T�i�i5a5`� 	 �_�R�[�oG ´s�o�kBp >qT>x�rH9B!�����~� <T��<]/���� U�@�y�d��������я��⏠`z�%�P
�M���]���n��� ��˟���ڟ����@I�4�m�X�����!Q�
V7.10b�eta1�V �@�p�@z=q�@��R�aʡC�  C5PB|ܣD7f@ �C�`���� D�� D�� C�`�`BY�䠃`C/�`p�R�r�`1�C�U�$�Bd�KNOW_M  ��U~VBdSV ��mi�-e :�ſ׿�z����
�PCσR�mAcMfc����8Plڢ	�Rܡ 3 �b�� ^�����S��ˠ`���I�iRL�MRfc�y�T�z��QCz����u8�J��6mSTfa1 1�V[
 0-e��$���  �ߙ߽߫��� ����4��)�;�M�� q�����������P��T�h�2s���NQ�<��a�3r�������l�4��������l�5"4Fl�A6_q��l�7����l�8�!�3l�MAD3V �^Vh�PARNUM  V[2πj�WSCH� ^U
�p� )@S%UPD����e\/�_CMPa_o�3PWPP'Wj�S_ER_CHK%|X�&/�+RS8�}�Ba_MO��/��%_�/\e_RES+_GrВv� ��n r?e?�?�?�?�?�?�? �?OO8O+O\OOO�_44q�><N?�O35�� �O�O�O53 �O�O _ 53^ _:_?_53� Z_ y_~_53� �_�_�_53�K�_�_�_52V 1�v�$1��@c����"THR_IN�R0"!W�(5dkfM�ASSxo Z�gM�Nwo�cMON_QUEUE �vը	6#0/��TNy U�!N�f�+�`END8�a?yEXE(u�> BE'p	�cOP�TIOw&;�`PR�OGRAM %��j%�`6o��bT�ASK_I�o~O?CFG ��o����DATArÖ.�@0�2��t� ��������g����� �(�ӏL�^�p���5��INFOr×Q�� �d=�ڟ����"�4� F�X�j�|�������į ֯�����0�B������Q� lI�� ?DIT ����>5�WERFLIx^c�i�RGADJ ����A�  ��?�#0�d�RG�a�}�y��?���Na�<@���ɖ%a�h�ϸ���2��5��`\hF]b2��2�A(d�t$���*��/�� **A:��#0����v��F�������W� Ab5�Ac	��-�?߬� c�u߇ߙ��߽����� N�I��)�;��_�q� ������������� �%�7�I�[�m���� ������������! �EWi{��� ��/��� Sew����� ��//+/U/O/a/ s/�/�/�/�/�/�/�/�??'?9?K?]?�? 	 ��?�?O�7��9O���OfOO�O����P?REF �%�Op�Op
۵IORI�TY�g��߱MPGDSP�qͿ�GU�g��ڶOG��_TGpʰ�r�j*RTOE�`�1��� (!�AFs`E�`s_~W�!tcp~_�]�!ud�_�^!�icm�_8o+QX�Yà���Oq)�� ��2oDoOp� ,omoPe\o�o�o�o�o �o�o�o�o;M4�qX��*)Sâ�MU�����?!�}�6��/���K��V��~ȁƺ�AG�,  ��@w���@����͏�E�t�C��O��Cղ߱PORT_WNUMS�����߱_CARTR�EP�@����SKS�TAW J�SA�VE ��	�2600H738B҈O�Or�`������LÉ7����7�Z�URGE_EN�Bʹ��aWF(�DOV{�EVWlPI�ձ�)�WRUP_DE?LAY ���=��R_HOT %��ֲ=�ɯZ�R_NORMAL��򲸯<�ܧSEMI��|Q���QSKIPȓ��� x}O��yO ��̿޿���=ϱ��� 4�F�X��|�jψϲ� ���Ϝ������0�B� �R�T�fߜ߮��߆� �������,�>��b� P����p��������(�2��$RB�TIF7_�ARCV�TM[BT�E�D�CRm��t� �Э�E8���E�d��C��B��\8������P(GŃ#���Añ��\7�´B������ ;��;����;�D�;��$;�< �Jl��Se  ����������	-?Q�GRD�IO_TYPE � ϝG]EFP�OS1 1���
 x?��Z@�< /�^��/v/a/�/ 5/�/Y/�/}/�/?�/ <?�/`?�/�??1?C? }?�?�?O�?&O�?JO �?GO�OO�O?O�OcO �O�O�O�O�OF_1_j_ _�_)_�_M_�_�_�_�o�_0o�_To��2 1����oJo��oFo�ojo�3 1��o�o�o�o`K�>S4 1�+�=w����S5 1��������u���,�S6 1� C�U�g����
�C���S7 1�؏����6�����؟V�S8 1�m����˟I�4��m��SMASK 1�z �������'XNOw������MOTEL�۫���_CFG ���b����PL_R�ANG�O�Q�OW_ER �����#�SM_DRYP_RG %�%������TART ��|�ʺUME_P�RO����&��_E�XEC_EN��zĄW�GSPD��pA�Iȓ�X�TDBd��v�RM��v�MT_ғ�Tw��E�OB�OT_ISOLC�خF�2�b���N�AME ���ÉOB_ORD_NUM ?|���H73�8 ~  �w��r����y�� �2�Dr�h��z��r� ���}�r����
r���x+��PC_T�IMEg�S�xE�S72320�1������LTEACH PENDANi�,,���7���P�Mainten�ance Con%s��$�"��T?KCL/Cٰp�����o� ?No Use��N�8��9���NPO��^����Y���C7H_L������	=��MAVA#ILSѸ�K������SPACE1 2�� �K�����2���K�L�b���?8�?�� ���IjAz�� �������': �_pW���� ���S'/:/ �_p/W/�/��� ��//#/?6?�/K? l?S?�?�/�/�/�/�/ �??1?3?�?GOhO?O QO�?�?�?�?�?�OO -O_}OC_d_v_]_�O �O�O�O�O�__)_o <o�_a_roYo�o�_�_ �_�_�oo%o8�o MnU��o�o�o�o �o�o�z�I�j� A��������� �/�!��E�f�x�O�a���2������͏ ߏ���%�4�U��j���r�����3��Ɵ؟ ����� �B�Q�r�5� ����������4ѯ� ����ǿ=�_�nϏ�@RϤ��Ϭ��ϥ�5�  ��$�6���Z�|ϋ߀��o��������ߥ�6 ��/�A�S��wߙ� ��������������7(�:�L�^�p���� ����������1��8E�W�i�{���; ������9 �N��G �e� E�
� �  e��� //%/7/g�V-� c�/+�/�d� � ��/??&?8?J?\? R/d/v.g:�?�;�?�/ �/^?O*O<ONO`OrO h?z?�?�?�?�O�O�? �?~O8_J_\_n_�_�_��O�O�O�O�O�_ `F @� +e�/ 9o_Ywa�Uo�o �o�_zj{o�o�o �oI[%/As �w����!�?� �'�i�{�E�O�a����Տ���\
Yo*���_MODE  e^@�S �e��_�Z�Uo~�П���	�� �CWOR�K_ADP�
^�dȡR  e�r g��Q�_INT�VALP���[�R_OPTION��� [��V_D�ATA_GRP �2��XpDPP ������C�1� g�U���y��������� ӿ	���-��Q�?�u� cυϫϙ��Ͻ����� ��'�)�;�q�_ߕ� �߹ߧ��������� 7�%�[�I��m��� ����������!��E� 3�U�{�i��������� ��������A/e S�w������W��$SAF_DO_PULS;��X��AZ�1!CAN�_TIMO�!U���BR �(�C��(�f0������Ē����S �����/ /�7/I/[/m//�/V���C,"2�$D��d�(�!�!�&�@�\
??.?*���)�/ ߠC4�w_ 3b  Tf��W?�?�?�?�9T D���?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_�����%_X_j_'Y�+a��Q;�o�*���p(]
�t� �Di�� -��,"���Q�� y�_o o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� �������� *�<�N�`�r���������̏-��T?���� +�=�O�a�s���ԏ�% ��ß՟�����/� A�S�X���-�0R2�S �U�]����ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ����� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�t�ߏ�ߪ߼��� ������(�:寧^� p����������� Y�����,".�@�R�d� v��������������� 	'9K]o� ������� #5GYk}��@������X�$_ �3/C/U/g/y/�/�/ �/�/�/�/�/	??-???Q?c?q:0/z?�?.�6�����?�=�	123456�78�R !B*�P
�8. �PO )O;OMO_OqO�O�O�O �A//�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_m�O$o6oHo Zolo~o�o�o�o�o�o��o�o 2DoBHU}���� �����1�C�U��g�y�����k;�j��ӏ���	��-� ?�Q�c�u���������0ϟ��
iD���%� 7�I�[�m�������� ǯٯ����!�3�E� oi�{�������ÿտ �����/�A�S�e� wωϛ�Z��������� ��+�=�O�a�s߅� �ߩ߻������߰�� '�9�K�]�o���� �����������#�5�G�$@d�v�[��������)"Cz � A�*   �(2�4A��A!+��0Ě22b�I�[m���0/���8��� !3EWi{�� �����//// �S/e/w/�/�/�/�/ �/�/�/??+?=?O?�a?s?�?�?�?�?�$�SCR_GRP �1�(ӈ�(ӿ� @�t ��
 �1 	 �3 AB 	D��"M�7GJO8O�qO��� nBD�` D��C�G�nK�R-20�00iB/165�F 567890�. �DX. R2�D7 �@B#
1�234�EAFnA� CV�1B&�3 �1�nAJBATY	ER�_�_�_�_�_~�\��H��0�TG�2&o5O6o\ono=FM/
Io�oEo��o���o��h,P�TpE  p�A�B���B�ff�B�33B�  �+v�5wAA��G # @
 _uA@�@oO  ?��wrH-p��JzAF@ F��`�r�=GC�  ��� ��D�/� h�S���w�7q_q�r��0����ʏ܄B��� 0��T�?�x�c�u��� ��ҟ�������*� �CZOH�m���  j�h��
�q@�r�O���=G��߯-p���@W\NCa�5�B$A�G��1Z��o�e �Y�
 {�����º���׸���Ŀ P��(!�'�9�K��1E�L_DEFAUL�T  XT���
 _�MI�POWERFL � ��w���WF�D n� w�^�R�VENT 1����`u���L!�DUM_EIP�M����j!AF�_INEk��B$!'FT��>��b�9!"o�� �Q߮��!RPC_MAIN�ߖ�������'VIS�ߕ	���F�o!TP9�PU=����d5��!
PM�ON_PROXY����e����Y�����f��*�!RDMO_SRV+���g��v�!R!T����h,e���!
��M�����i��!RLSgYNC5	8��>Z!ROS�ρ��4I�!
CE>[�MTCOM����k��!	�CONS���l�>u� b9�/A��w� ���/�@///�+/�/O/a/Q�RVI�CE_KL ?%��� (%SVCPRG1�/:�%2??� 3+?0?� 4S?X?� 5{?�?� 6�?�?� 7�?�?� HTO<9O K�$ ��HO�!�/pO�!?�O �!E?�O�!m?�O�!�? _�!�?8_�!�?`_�! O�_�!5O�_1^O�_ 1�O o1�O(o1�O Po1�Oxo1&_�o1 N_�o1v_�o1�_ 1�_@B1�_�/�"�  �/� ��1��� ��@�+�d�O����� �������͏��*� �<�`�K���o����� ̟�����&��J� 5�n�Y���}���ȯ�� �ׯ���4��X�j� U���y�����ֿ�������0��Tϖz_D�EV ����MC:\� 
�]n�OUT`�h���j�REC 1Ÿ�uh��� �� 	 \������؁3�lu:��c�n�
� �Tpvj6� sS��  �����  �  Пл�u��X�Wr 1��h�=h�Y��ů� ����h�U+h���2���� �����'�M�;�q�_� ������������ �#�I�7�m�O�a��� ����������! E3UWi��� ����A/ QwY����� ��/+//O/=/s/ a/�/�/�/�/�/�/�/ �/'??K?9?o?�?c? �?�?�?�?�?�?�?#O ���O)OOQO�OuO �O�O�O�O�O_�O)_ _9_;_M_�_e_�_�_ �_�_�_o�_%o7oo [oIoomo�o�o�o�o �o�o�o3!WE {�o����� ��/�A�#�e�S��� w��������ŏ��� �=�+�a�O�����y� ����ߟ͟���9� �I�K�]���������xۯ�׽�V 1���� (ӯ&���TOP�10 1���
 ��,�v�����@��YPE��l�HEL�L_CFG ��{�h�	�  x��B�RSR� �/�h�Sό�wϰϛ� �Ͽ���
���.��R߰=�v߈ߚ������%�����ߨ�������������װ�2h�d����϶�HK 1�ݻ 
��������� ������+�=�f�a� s�����������h�϶?OMM �ݿ�βFTOV_EN�B���ƺOW_R�EG_UI=ͲI_MWAIT:��.mOUT^�o	wTIM^����VAL~p_UNcIT9�ƹLCW WTRY^Ƶ���MON_ALIA�S ?e	�he�Vhz���� R���/�%/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?�/ i?{?�?�?J?�?�?�? �?O�?/OAOSOeOwO "O�O�O�O�O�O�O_ _+_=_O_�Os_�_�_ �_T_�_�_�_oo�_ 9oKo]ooo�o,o�o�o �o�o�o�o#5G �oX}���^� �����C�U�g� y���6�����ӏ��� ���-�?�Q���u��� ������h����� )�ԟM�_�q�����@� ��˯ݯﯚ� �%�7� I�[���������ǿ r�����!�3�޿W� i�{ύϟ�J������� �Ϥ��/�A�S�e�� �ߛ߭߿���|���� �+�=���a�s��� B�����������'� 9�K�]�o�������� ��������#5G ��k}��L�� ���1CUg�y#�$SMON�_DEFPRO ������ *S�YSTEM*  �ȏRECALL� ?}� ( ��}.xcopy� fra:\*.�* virt:\tmpback��=>portuc:18700 !`/&/8/J/#}2��s:orderf?il.dat�,��/�/�/�/]!)�mdb:�,�/?/?�A?T*-���0  ?�?�?�?X&�r?/�O(O:OLO }x�yzrate 11L�?O�O�O�OU)�9�$:manut�entionpi�nceauto.;tp�5emp�/_/_A_TOfA6kM�O_ �_�_�_U_gOy_�_o(.o@oS+0�On�_ ? o�o�oOo�O�O|o�o (:L__�_� ���_o��$�6� H�[�������Ə Y/k/�/�C��&�8�J� �/���o�����ȟ[? �??��"�4�F��?� ���C�����ʯ]ooo ����$�6�H�ۏ�v� ������ƿY�m�}���  �2�D�ן�|���� ����U�g�xϋ��.� @�S�e��N߬߾� ѿ�~�ϙ�*�<��� a��υ�������� p�ߕ�&�8�J�ݯ�@��������[�/b�ouvre�bu������$6H[�*b�prog1���?� ��[�m����"4 F��������� W�i����/0/B/�� �����/�/�/�� n	�/,?>?Qc�/ �?�?�?O?�t// �?(O:OLO_/�?�/O �O�O�O�/�/x?�O$_ 6_H_[?m??_�_�_��_�d�$SNPX�_ASG 1������Q�� P� '%�R[1]@1.Y1�_i?��c%o Do'ohoKo]o�o�o�o �o�o�o�o�o.8 dG�k}��� �����N�1�X� ��g�������ޏ��� ���8��-�n�Q�x� ����ȟ�������� 4��X�;�M���q��� į���˯ݯ��(� T�7�x�[�m������� �ǿ����>�!�H� t�WϘ�{ύ��ϱ��� ���(���^�A�h� ��w߸ߛ߭������� $��H�+�=�~�a�� ������������ D�'�h�K�]������� ����������.8 dG�k}��� ���N1X �g������ /�8//-/n/Q/x/ �/�/�/�/�/�/�/? 4??X?;?M?�?q?�? �?�?�?�?�?OO(O TO7OxO[OmO�O�O�O��O�D�TPARAM� ��U�Q ��	��JPXT�XP�XOFT_K�B_CFG  �%S�U?TPIN_S_IM  �[4V��_�_�_7P�PRVQSTP_DSBn^�4R�_"X�@SR ��qY � &� �_/o%P<VT�HI_CHANG�E  %T�\WOaGRPNUM�OV djOP_ON_ERRYhZY�a?PTN qUc`�AKbRI�NG_PRy`�n��@VDTsa 1�<Ya`  	8W"X 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� a�^�p���������ʟ ܟ� �'�$�6�H�Z� l�~�������Ư�� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�y�vψϚ� �Ͼ���������?� <�N�`�r߄ߖߨߺ� �������&�8�J� \�n���������� �����"�4�F�X�j� ���������������� 0WTfx� ������ ,>Pbt������?SVPRG�_COUNTOVq��a^U"ENB�o�	%M3#|eA/UPD� 1�kT  
�%R�/�/�/�/�/ �/�/??,?>?g?b? t?�?�?�?�?�?�?�? OO?O:OLO^O�O�O �O�O�O�O�O�O__ $_6___Z_l_~_�_�_ �_�_�_�_�_o7o2o DoVoozo�o�o�o�o �o�o
.WR dv������ ��/�*�<�N�w�r� ��������̏ޏ�� �&�O�J�\�n����� ����ߟڟ���'�"��4� +YSDEBU)G y �J�da)l�SP_PASS%�B?~�LOG [�x%c#J�9G�T�  �]!J�?
MC:\��Z���_MPC��x%,�$>�x!�\� x!��SAV ѳ��Ф�J��SV�_�TEM_TIM�E 1�x)��(�Ѡ^ͤ]ȯ)T1?SVGUNSs %�'a%�	�ASK_OPTION �x%]!'!)�_DI���4/E�BCCFGg �л�� ���ό�`������� �������7�"�[�F� �jߣߵߠ������� ��!��E�0�B�{�f� ������������J�	�8�
�k�}��� Z�����������c� ;���#I7m[� ������ 3!WE{i�� �����//-/ //A/w/](H��/�/�/ �/�/]/?�/?9?'? ]?o?�?O?�?�?�?�? �?�?�?�?OGO5OkO YO�O}O�O�O�O�O�O _�O1__U_C_e_g_ y_�_�_�_�/�_�_o -o?o�_coQoso�o�o �o�o�o�o�o) M;]_q��� �����#�I�7� m�[��������ŏǏ ُ���3��_K�]�{� �����ß��ӟ��� �/�A��e�S���w� ��������ѯ���+� �O�=�s�a������� Ϳ���߿��%�'� 9�o�]ϓ�I��Ͻ��� ����}�#��3�Y�G� }ߏߡ�o��߳����� �����1�g�U�� y���������	��� -��Q�?�u�c����� ����������; M_���q��� ���%I7 m[}���� �/�3/!/C/i/W/ �/{/�/�/�/�/�/�/ �//??S?	k?}?�? �?�?=?�?�?�?OO =OOOaO/O�OsO�O�O �O�O�O�O�O'__K_ 9_o_]_�_�_�_�_�_ �_�_o�_5o#oEoGo Yo�o}o�oi?�o�o�o �oC1Syg���v�p�$TBC�SG_GRP 2�Շu� � �q 
 ?�  ���� �@�*�<�v�`�������r�s��|d0�ہ?�q	 H�D)̪�&ff�����B\�r�!�N�333?���!�#��L�͇�L���ޱ�C�����ϖ��CA�CA4����Ř@�� �����Ř���HA���@ �p������¯�����
�կ�5�R�a�7�p�  ,	V3�.00�r	r2;d7a�	*������r��k���(�p7� q㰵��  ������M�&�-ÿqJ�CFG هu��q�-��W�r��-ς���� �϶ʐp������ ��� $��H�3�l�W�iߢ� ���߱��������� D�/�h�S��w��� �����
���.��R� d��r�`o�����=��� �������� D/ hz��Y��� ���q�A�Q Se������ /�/=/+/a/O/�/ s/�/�/�/�/�/?�/ '??K?9?o?]??�? �?�?�?�?�?�oO)O �?IOkOYO�O}O�O�O �O�O�O__1_�OA_ C_U_�_y_�_�_�_�_ �_	o�_-oo=o?oQo �ouo�o�o�o�o�o�o )M;q_� �������� 7�%�[�I�k���;O�� ��͏w������!� W�E�{�i�����ß՟ �������-�S�e� w�1�������ѯ���� ���)�+�=�s�a� ��������߿Ϳ�� �9�'�]�Kρ�oϑ� �ϥ���������#�5� ߏM�_��ߡߏ��� �����������C�U� g�%�w�������� ��	����?�-�c�Q� s������������� ��)_M�q ������% I7m[}� �A���/�3/!/ C/i/W/�/{/�/�/�/ �/�/?�//??S?A? c?�?�?�?g?y?�?�? O�?+OOOO=O_O�O sO�O�O�O�O�O�O_ __K_9_o_]_�_�_ �_�_�_�_�_o�_5o #oYoko/�o�o/Qo �o�o�o�o/U Cy��[m�� ���-�?�Q��u� c�������Ϗ���� ��;�)�K�q�_��� ������ݟ˟��� 7�%�[�I��m����� ��ٯǯ��wo�o'�9� ��W�i�����ÿ�� �տ��/�A���e� S�u�wωϿ������� ����=�+�a�O�q� s߅߻ߩ�������� '��7�]�K��o�� �����������#�� G�5�k�Y�����K��� ��������1A CU�y������	�-Q; s w{ {��{�$TBJO�P_GRP 2��C� / ?�{	���ܵ�K�� `p�p� ��� � � �{ @w�	� �D)�+%C2
C랔{��G"333O!>̓��K/! LY p$<���d+!? !p$B�`  A�A$�����'+/=/O%O"�/��*<+�~-C/  B�{@!/?��/�/F'p%�%p=�=��5<ҙ*"P!p!�Cz!0�$�?�;�C�6���C�p��.�?K�%�p ;��:CA�i��"P$C�C4�?�VO�?�?m(�Oj;(A�S=�/JhAH�0 YO��OiO{O_+^fff?U<:f�/F !�0 ?B�@f_x_+_�_�Y�_ �_�_�_o�_�_!o;o %o3oao�omo'o�o�o �o�o�o"�D�{� � �G%	V3.�00�r2d7�*mp�v{�w GO �~�d� G�0G��� G�| G�:� G�� G��� G�t G�2� G�� Gݮ� G�l G�*� G�� HSޖrFj` �~�� F�q � G�X G/� GG�8 G^� Gv� G�ĺs�4� G�� G��� G�\ G�{ =p =#�
|8(1Cq�j�k�}�5{��?�X�����ESTPARb�po��HRրABLE 1ݵI��{���� ��v�������z�*��	��
������{������N�RDI����@!�3�E�W�i�єOٟ������+�=��Sן� �����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� �֠گ	���~����� ��`�r����������~{�NUM  C�� � ��̐�_CFG ��d��!@�IMEBF_TT܁pս逦�VERʓ�������R 1ߞ� 8x{dv� F��  � �%�7�I�[�m��� ������������!� 3�E���i�{����������������_b̐/� �  kX����T��6���9��I���/ �LTA_ż6���L�:6���B���� 7�����/ 
��:���);^�g]o  ŋR�ƙs/ �Vdà��/ �W����
�/� [X�s%��	/���_^���@���ӀMI_CH�AN�� �� �#D_BGLVL�����ҁ� ETHERA�D ?��� ��������/?ˈ� oROUT��!���!54S?&<SNM�ASK�(���!255.�5Ys�?�?�?�YsӀOOLOFS�_DI�pM%�)O�RQCTRL I��ɖ���1NT O UOgOyO�O�O�O�O�O �O�O	__-_?_Q_c_�u_�\O�_�_�_ЃPE_DETAI�(��:PGL_CON?FIG �d�t����/cell�/$CID$/grp1�_FoXojo|o�oD��?�o�o�o�o �o7I[m � ������ ��E�W�i�{����� .�ÏՏ������� A�S�e�w�����*�<��џ�����+���} ��a�s���������)��_�­����*�<� N�`�r���������̿ ޿���&�8�J�\� nπ�Ϥ϶������� �ύ�"�4�F�X�j�|� ߠ߲���������� ��0�B�T�f�x��� �������������,� >�P�b�t�����'��� ��������:L ^p��#����� $`�E�User Vie�w 4oXjI�}1�234567890�������X@ c/��;2q =/O/J�s/�/�/�/�/ �/=�//C3�/!? 3?b/W?i?{?�?�?�?�/�/<4�?OOF? ;OMO_OqO�O�O�?�?<5�O�O�O*O_1_�C_U_g_y_�O�O<6 �_�_�__oo'o9o Ko]o�_�_<7eo�o �o�_�o�o/Apo�o<8I���o �����%�TF�� �ECameraFx���������ҏ�����E ��9�K����x����� ����ҟ�`�+/�'� ��K�]�o�������� ɯۯ�8��#�5�G� Y�k�2�pu`�?��ÿ ������/�Aϸ� e�wω�Կ�Ͽ����� ���~����?M�_ߞ� �ߕߧ߹�����T�� �%�p�I�[�m��� ��ߐ��O����:�� 1�C�U�g�y��ߝ��� �������	-? ��_������ ����9K] �������R ���o!/3/rW/i/{/ �/�/�/(�/�/�/D/ ?/?A?S?e?w?��� ��?�??�?OO)O ;OMO�/qO�O�O�?�O��O�O�O__�?��9 !_Z_l_�O�_�_�_�_ �_�_aOo o2o}_Vo�hozo�o�o�o'_qt	a�0�o�o	Ho-? Qcu��_��� ���)�;�M��o�l1Y������ɏۏ ����#��G�Y�k� ��������şן�`��l2��/�A���e�w� ��������6����� R�+�=�O�a�s������l3��˿ݿ��� %�7�I�[�үϑϣ� ����������!ߘ��l4-�g�y߸ϝ߯� ��������n��-�?� ��c�u�����4��l5����T�9�K� ]�o�����
������ &���#5GY���l6e������ �/��Sew �������lz  w	+/=/ O/a/s/�/�/�/�/�/<�/�+   /	/ '?9?K?]?o?�?�?�? �?�?�?�?�?O#O5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_ g_y_�_�_�_�_�_�_ �_	oo-o?oQoco�,�  
s (  }� ( 	 so �o�o�o�o�o�o %'9o]���:}j: �K� � ��D�V�h�z��� ��u�ȏڏ�3�� "�4�F�X�j������� ����֟�����0� w�T�f�x��������� ү���=�O�,�>�P� ��t���������ο� ���]�:�L�^�p� �ϔ�ۿ������#� � �$�6�H�Zߡϳϐ� �ߴ���������� � 2�y�V�h�z��ߞ�� ��������?��.�@� ��d�v���������� ���_�<N` r�������% &8J\�� �������/ "/i{X/j/|/��/ �/�/�/�/�/A/?0? B?�/f?x?�?�?�?�? ?�?�?OO?,O>OPO�bOtO�O�?�p@  �B�O�O�O�C�G�`����O_&_8_J_ \_n_�_�_�_�_�_�_ �]_o o2oDoVoho zo�o�o�o�o�o�o�_ 
.@Rdv� ������o�� *�<�N�`�r������� ��̏ޏ���&�8� J�\�n���������ȟ ڟ����"�4�F�X� j�|�������į֯� ����0�B�T�f�x� ��������ҿ���� �,�>�P�b�tφϘ�Ъϼ����I(A ��O�$TPGL�_OUTPUT ���1�1 ���,�>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p���������������  2345678901����%� 7�I�Q��2��x����� ������j���,>P��}Z��� ��bt $6 HZ�h���� �p�/ /2/D/V/ � /�/�/�/�/�/�/ ~/�/?.?@?R?d?�/ r?�?�?�?�?�?z?�? O*O<ONO`OrO
O�O �O�O�O�O�O�O�O&_ 8_J_\_n___�_�_ �_�_�_�_�_o4oFo Xojo|oo�o�o�o�o�o�o�o��}��0B Tfx��}@�Ͽ������( 	  ����*��N�<�r� `�������̏����ޏ ��8�&�H�n�\��� ������ڟȟ�����4�"�X���OFF�_LIM#��������t�N_�SVx�  �����P_MON ��َ��������S�TRTCHK ��Պ�-��VT?COMPAT��)����VWVAR �뿭"�N��� R � d���Ң��_DEFPROG� %�%
OU�VREPINCE{  ��AUTO{�~��ISPLAY#���INST_M�SK  � ~кINUSER��ִLCK(��QU?ICKMENL�ִoSCREk��~*�tpscִ�(����Ɋ���_��S�T���RACE_�CFG ��jL�Ϡ	��
?��~��HNL 2�L��S� y�?�Q� c�u߇ߙ߽߫�����ITEM 2�+۟ �%$� � =<�B�T�\� G !b�j�v�&� ����4����j� ����i������� ��@�0�B�T�n�x��� ��Hn���� ,�P�"4�@ ���d��� L�p�K/�f/� �/�/ /�/$/v/�/Z/ ?~/*?P?b?�/n?�/ �/?�?2?�?OOz? :O�?�?�?FO^O�?�O �O.O�OROdO-_�OH_ �Ol_~_�O�___�_ <_�_`_o2o�_�_�_ �_�_�_joo�o�o�o \o�o�o�o�ot ���4FX� *��N�`��l��� Ï�ޏB���x�*� ���w�ҏ������ȟ ڟ>��b�t��� ��� V�|���򟲯�(�:� ��֯p�0�B���N�ʯ ܯ�� ���$����Z���~���Y���S���|��^��  ���^� ѵ���
 ��������d�R_�GRP 1���� 	 @�� L�^�H�~�lߢߐ����ޠ���������%�x�I�4�?�  d� v�`��������� �����8�&�\�J���`n���������	,���� )�SCB 2�z� O�L^ p������d��X_SCREEN� 1�7�
 �}�ipnl/g?en.htm�<�N`r�&�P�anel setup�}������/"/ ��Z/ l/~/�/�/�/+/�/O/ �/? ?2?D?V?�/�/ �?�?�?�?�?�?]?�? �?.O@OROdOvO�O�? �O#O�O�O�O__*_ �O�O`_r_�_�_�_�_ 1___U_oo&o8oJo \o�_�o�_�o�o�o�o��o�ouo�UALR�M_MSG ?7���� _zQ c������� ��6�)�Z�M�~�2u�SEV  @}i��0rEt��z������A��   B������7��%� 7�I�[�m���������ǟ՗��1��Ƌ �?�4����A��*SYSTEM*&��V8.1079 �G�1/30/2013 A 7���5�"�UI_ME�NHIS_T �  8 $q�T__HEAD��}�ENTRY ���$DUMMY2�  ��3�� � j�OUSEt����$ACTIO�N��$BUTT�ˤROW͢COL{UṂTIME���$RESERV�ED��j�PAN�EDATt� �� $PAGEU�RL }$F�RA�)$H�ELP�PA'�TER1+�<���H����H�4F�5F�6F�7�F�8+�INB�VAx ���	�STAT*�⥥1r����� �j�USRVIE�Wt� <Ġn�Uz!��NFIG���FOCUS��PR�IM!�m�����T�RIPL*�m�U�NDO_t�t� � $4�ENB~��$WARNJ�|����_INFOt��y��_PROG� %$TAS�K_I��t�OSIKDX��R��`��TOOLt� 4o $X��$��r��Z��ߡ$P��R�°�NU�9`�	U&�t��������9E��`�OFF��u�� D{���O?� G1��)�Q����GUN_WIDT�H  ��K�_�SUB��  
F`�RT���t�	���$D����OR�N��RAUX��T���ENAB-���V�CCM��� �
$VISʠ_TkYPɳC(�RA��GPORTХ�A�C�z��N(�%$EX��)_��$��_F�P�ʣ�P� A��a�LU� �$OUTPU�T_BM��ӝ��MR_���h ����+��DRIV����SE�T_VTC���B�UG_CODɴM�Y_UBYȴ6�	 ����ʠE��,���:��f�x�O�HANDE1Y��E�8pULX�P���AL_���GD_SPACIN���RGT�������0�����U�RE����U��w� �������  ��RG���PNT�CR\���� dġXr��FLA���	T�A�XS���SW��_)A��y���S��O��BA��zy�	$E��UE���y�Ҁ��+HK�� �
зMAXvER��MwEAN�	WOR���z-MRCV��� ��ORG9pT_C&P )�
REF���- �i ��яN��b b1��_RC���� 8���M���M�ր��� �P�űG]�����$GROU�P����:&�� ���2p C�REǰw��$��Ab"N!HK��S�ULT���CO�VE����a NT6��%���&���&ձ�#m L6��%F��%����'ձ���9��0 &z#PA�u� z#CACHO�LOV*4@1��E9����C_LIMmIf3FRn8TDn8N�$HO��=�.0�COM������OB�O�8(� �!$IN�_VP�����2_S�Z3�#�56�#�51�2���8R��:TKQ��8o0�8WA5MP�BJFAIo0G��?0ADrIU�IMRyE $�B_SIZ/$�PM��ND� P�A�SYNBUFP�V�RTD�E�D�A�3O?LE_2D_��EmW�PC��TUq��@0Q� �EECCU��VEM��)54Ro6� ��$��� C�KLASv�	�V�LEXE5G���� �z!O�FLD6d�DE�CFI�@�W�� �W-;�s� (����
��QǠ�ѡ ��_��L�#���8 hP �1���!��K�$��$�=�E�!}�C�U�%$"A7
�@PS�Kt4M:&�e  ���TRbUt�� $p TIT-���A0=�OPɤ��VSHIF:��`��|!#����URO�d _R�@�+t H�C=u��L�^�p�o0`���qi �ҏsTI�!N�tSCO'r�sC�� ��S¨�SwS£vS� �wS¾x����Ꞣ���s�ED���w� m SM7�A��$ADJ�`K�%�UA_{"u�A��g�}�LIN.����ZABC������
�QZMPCF���  C��J���LN�`�a��I��� ���1� ���CMCM��C�3COART_6��Pa? $JT�N�D�1Z�k�d���p���ΎUXW����UX!E�񞖙�_���u����������ɖ!ZP�5��r�������Y:��Dc� y�2v�/�IGH���h?�(p ���$ � � �d7ۀ$%Bm KK�]a_�b�#u�RVn0F��cOVC��O�D��$�`(��Ǳǡ
�Iݣ�5}D�TRACEJ��V�R��SPHER>�� ! ,p 1��G�Y��$�DEF~x�?%���c���^�(%�ހx���t�����ѿ �������*�O�:�`s�^ϗϢ�T�IN���  c��Ϧ�_�T`H��1 c���(�� ���(/SOFT�͡/GEN��K?�current=�menupage?,153,1��T�8f�xߊ߀� �.�962A���������߭߿�36��Z�l� ~����������� ����7�I�[�m�� �� ����������� ��3EWi{�� .����'��ѶSew� ������// +/�O/a/s/�/�/�/ 8/J/�/�/??'?9? �/]?o?�?�?�?�?F? �?�?�?O#O5O�?�? kO}O�O�O�O�OTO�O �O__1_C_.@y_ �_�_�_�_�_�O�_	o o-o?oQo�_uo�o�o �o�o�o�opo) ;M_�o���� ��l��%�7�I� [�m��������Ǐُ �z��!�3�E�W�i� T_f_����ß՟��� ���/�A�S�e�w�� ������ѯ������ +�=�O�a�s������ ��Ϳ߿�ϒ�'�9� K�]�oρϓ�"Ϸ��� ������ߠ�5�G�Y� k�}ߏ�z��������� ����"�C�U�g�y� ���,�>�������	� �-���Q�c�u����� ��:�������) ����_q���� H��%7��[m��������$UI_PAN�EDATA 1�����  	�}��/ /2/D/V/h/ ) j/�/�$��/�/�/�/ ??z/7??[?m?T? �?x?�?�?�?�?�?O��?3OEO,OiOvI� ���B�/�O�O�O �O�O _SO$_�/6_Z_ l_~_�_�_�__�_�_ �_�_o2ooVo=ozo �oso�o�o�o�o�o
}L+v�H_M_q ����o�>_�� �%�7�I��m��f� ����Ǐُ�����!� �E�W�>�{�b����� $6�����/�A� ��e����������ѯ ���\�� �=�$�a� s�Z���~���Ϳ��� ؿ�'��KϾ�П�� �ϥϷ�����.���� ��5�G�Y�k�}ߏ��� �ߚ����������1� C�*�g�N������ ����X�j�(�-�?�Q� c�u����������� ��)��M_F �j����� �%7[B� ������/!/ tE/��i/{/�/�/�/ �/�/</�/�/??A? S?:?w?^?�?�?�?�? �?�?O�?+O��aO sO�O�O�O�OO�O�O d/_'_9_K_]_o_�O �_z_�_�_�_�_�_o #o
oGo.oko}odo�o0�o�o8OJO}��o !3EWi)�o� U}������ {8��\�C�U���y� ����ڏ�ӏ���4��F�-�j�v�TCNK�$�UI_POSTY�PE  TE� 	 v��͟��QUICKM_EN  �����П��RESTOR�E 1TE  �]�G�A�S�w�mr����� ��ѯ㯆���+�=� O��s���������f� ȿڿ�^�'�9�K�]� o�ϓϥϷ������� ���#�5�G�Y��f� xߊ������������ ��1�C�U�g�y��� ��������ߚ��� ��:�c�u�������N� ��������;M _q�.����& �%7�[m ���X���x/!/ۗSCRE��?�u1�sc<�u2\$3�\$4\$5\$6\$7�\$8\!��USER�> C/U"T= ^#ksTf#�$4�$5�$6�$�7�$8�!��NDO_CFG ����`�a��PDATE� �)�N�oneޒ� _IN/FO 1�&Q0��0%'/l?x8Z?�?~? �?�?�?�?O�?+OO OOaODO�O�OzO�OԜ�>1OFFSET ��OS5�� __0_B_o_f_x_�_ �_�_�O�_�_�_o5o ,o>okoboto�o�[ ���m
�o�o�HUFR�AME  �d�6;1RTOL_A�BRT932rEN�B;,xGRP 1�	0���Cz  A��s�q�a������v��*z��U[x1J{MSK � ^uQ3LyNq�%I:%�o��ݒVC�CM_PAp �
<%~VSCAM1 *ߏ�焣����5��V��MRwr2��ҀI�?��	с��	ֆ��Z�1B��5�A�@�pp�pȣ� 	�o����������<������uA����T�Z� B���o�Z�s� ����۟����ܯǯ � �$��!�Z���;����{���ƿy������I�SIONTMOU4:p^�˅���"�f`��f`��@�q FRk:\�\0A\�� �� MC�T�LOGa�   oUD1T�EX�����' B@ �������ϙ������ � � =	 1- �n6  -��� t������, ֌�_�=����h����z�TR�AIN��$�4��� (��h��ݧ� ���������"�4�j� X�n�|�����﯆/LEXE<��1�1-80��MPHA�SE  &53�k���R 2�
 ��]�o��������a������  ���� $6*1l����������� ��s����������G	no�pqrs�tuvw Z�~��� ����./f</ n`/r/��/�/�/�/�//h$/?H/&? L?~/p?�?�?�?�?�? /? O2?$O6Oh?ZO�lO~O�O�OD�{u�3��? �OO__LO>_P_b_�t_�_D��D	��BH
�O�_�O�_ o4_&o8oJo\onoH��@~		�3�
�
��Æ�o�_ �o�oo&8J�|o�3�
�
ghijk�@ \��o��o�o����&�8�ƃ��SHI�FTMENU 1,>�c�<��%�ϖ�&���t���ӏ���� 	����?��(�N��� ^�p��������ʟܟ �;��$�q�H�Z����~�T��[�K��	VSFT1��~VSCAM�S�5ذ?��!�@`��G�  A�ٰ8*ٰٰ��p*�$����"�!����9�L�̦MEP �a�/� T�MO����zR�WAIT?DINEND � �|w���OK  O�ȵ��ԿS迻�TI]M����G�� 5�ǿX��8��8�%���RELE9�h�s�f��TM��s����?_ACTIV��1����_DATA 	[�2�%��h�,���RDISg�����$ZABC_GR�P 1۩I�,�qp�2p�t�ZMP?CF_G 1�v��I�0�������MP¨�۩/��'��8��'�s�8����0��_����?����� ���/����V�������`�[������@�������Ѕ������P_CYLIN�DER 2��� Н� ,(  *m~��j���� ��% gH�lSe�� ���-/��D/ +/h/O/��/�/��=�s2 ۧ4� �� �/<�~�3??W?e:h�/�?�7��1A�;�SPHERE 2!M�/�?R/�?O �?8O�/�?nO�O��O CO)O�O�O�O�OWO4_ F_�O�O|_�O�_�_�_��__�_oo��ZZ�� ���