��   D�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A 
  ����CELLSET�_T   �w$GI_STY�SEL_P }7T  7ISO:iRibDiTRA�R�>�I_INI; �����bU9AR�TaRSRPNS�1Q234�5678�Q
TROBQACKSNO� �)�7�E�S �a�o�zU2 3 4 5 6 7 8awn&GINm'D�&��) %��)4%��)P%�̖)l%SN�{(OU���!7� OPTNAA�73�73.:B<;�}a6.:C<;CK;C�aI_DECSN�A�3R�3�TRY�1��4��4�PTHCN�8D�D�INCYC@HG��KD�TASKOK �{D�{D�7:�E� U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V�8�Tb@SEGq�Tp��T�@REQ� d�drG�:Mf�GJO_HFAUL�Xpd�dvgALE�  �g�c�g�cvgE� �H<�dvgNDBR�H�dgRGAB�Xtb�� �CLML�Iy@   �$TYPESI�NDEXS�$$�CLASS  O���lq�����apVIRTUA�Li{q'61ION�  ��c��q�t+ UP0 ��u�qSty�le Select 	  ��r�u�Req. /Ec�ho���yAck����sInitGiat�p�r�s�t�@�O�a�p���	���  ����*�������q��������q��sOpt�ion bit �A��B����C��Decis�c�od;��zTryo�ut mL��Pa�th segJ�n�tin.�II�y�c:��Task �OK��!�Manu�al opt.r��pAԖBޟԖC��� decsn �ِ�Robot interlo�|"�>� isol3���C��i/�"�z�ment��z�ِ�����_�status��	MH Fau�lt:��ߧAle�r��%��p@r 1�z L��[�m��+�; LE_COM�NT ?�y�   ��䆳�Ŀֿ �����0�B�T�g� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼�����������U������  � ��ENAB  ���u���������ꐵMENU�>�y��NAME {?%��(%$*4� ��D��p2�k�V���z� ������������1 U@Rdv�� �����* <u`����� ���/;/&/_/J/ f/n/�/�/�/�/�/? �/%??"?4?F?X?j? �?�?�?�?�?�?�?�=