��   to�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����UI_CONF�IG_T  �$ 5$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY5]0�ODE�
1CWFOCA �2C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� �4 TOUCH�P{ROOMMO#{?$4 ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"��%�!BA�!j ?��"BG�%$PM��X_PKT�"I�HELP� MERޱBLNK$=EN�AB�!? SIPMoANUA� &�USTOM0 �t $} RT_OSPID�p4Cx4n*PAG� ?^�DEVICE�9S�CREuEF����7N�@$FLA�G�@ [2�1 � h 	$PWD?_ACCES� E �8�C�!�%�)$LABE� '	$Tz j�0q!�@D�	�3USRV�I 1  < �`� vB�wAPRI�m� U1�@�TRIP�"m�$�$CLA�0 �����A��R��R�@VIRTT1�O�@�'2 )�7)��@�R	 ,��)?���RPS�SQ�� , ��Y03_��
 ���Aw_�_�_�_�_�_�_ s_oo,o>o Pobo�_�o�o�o�o�o �ooo(:L^ p�o������ }�$�6�H�Z�l�� ������Ə؏�����  �2�D�V�h�z�	��� ��ԟ������.��@�R�d�v���PTPTX���|���� s Ǖ����$/soft�part/gen�link?hel�p=/md/tpmenu.dg�� $�6�H�Z��&��pwd�����˿ݿ ���%�7�I�[�� ϑϣϵ�����h�zπ�!�3�E�W�i�?T���AMV/VS��($�ϻ������������AQ,�._��8����ߜ�lS��NQd��P���  ��X��Z@����f���8*��Ca2 1�EP�R \ }|Y0REG �VED�����w�holemod.�htm"�sing}l3�doubJ��tripb�?brows{�f� ������������/Aj�����/�d/ev.s8�l�]�� 1�	t���� e�5GY#}�p����� �@ //*/</N/`/r/�/ �/�/�&�0/�/�/�/ ? ?2?5����e? w?�?�?�?�?�?�?�? OO+O=OOOaOsO�O �O�Ow�O�O�O�O_ _1_C_U_g_y_�_�_ �_�_�_�_�_	oo-o �hozo�o�o�o�o�o �o�o
?.@! v�??Q?7o��� ���%�7�`�[�m� �������Ǐ����� �O��E�W�i�{��� ����ß՟����� /�A�S�e�w���Woį ֯�����0�B�T� f�a����k�}�ҿ� ����,�'�9�K�t� oρϓϼϷ������ ���#�L�G�Y�'�y� sߡ߳���������� �1�C�U�g�y��� �������ﳯ �2�D� V�h�z����������� ��������.@��	� �������� �%7`[m �������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?�|?�?�?�?�? �?�?�?OOBOTO�#O5O�O�O�J�$U�I_TOPMEN�U 1u@�A�R 
X��AT1)*def�ault_?H=	�*level0 *P �O�5_�4_F_�tpio�[23]�tpst[1yXoP�O�_�Z_S_�_�_�_�	�menu5.gi5f�
*a13/i(c�1/k)b4/ko�Q��{o�o�o�o�o�o�o S2�o%7I[m ��������!�3�E�W�i�{�����prim=*ac?lass,5��Ï�Տ�������13�H�Z�l�~�������page,153,1��Ο���(�����8��O� a�s��������ͯ߯���L9�@�A�O M�]?��Q=�wo��V�ty�]r_�Qmf[�0�_�\	��c[1364yW�59yX�Qeo��A�#h2Wo-m�� CjOo9gVj�ϊd-�?� ��0�B�T߫�xߊ� �߮�����a����� ,�>�P��ߡ�2b�� �������n﬏�'� 9�K�]�����6����� ����������1��$�6HZl����ainediE�������zwintp���(:L^p O6�A8�z��V�_H� ���//,/>/P/ �_p/n/�/�/�/�/�/ �/?)?�oM?_?q?�? �?�?���?�?�?OO %O�?IO[OmOO�O�O �ODO�O�O�O_!_3_ �OW_i_{_�_�_�_@_ �_�_�_oo/oAo�_ eowo�o�o�o�oNo�o �o+=�oas@�������5� �Y�k���u�#?5�ӺAs��R�w�ſ_�u�� *�,φ�����Æ��h.�|�R�6_�u7�� ���Ϸ�ɟ۟���V #�5�G�Y�k�}�������ůׯ��������1	�G�Y�k�}��� ����ſ׿���Ϝ� 1�C�U�g�yϋϝ��� ��������	�ߪϼ�6"�W�i�{ߍߟ�����74��������� #�G�Y��/@��� �����������z� �B�T�f�x������� ��6?��	-?Q �u������ p);M_� ������l/ /%/7/I/[/m/��/ �/�/�/�/�/z/?!? 3?E?W?i?�/�?�?�? �?�?�?�?�?O/OAO SOeOwO2�D�Oh�2� ���O�O__=_<_N_ `_�Ol_�_�_�_�_�_ �_oo��Ko]ooo�o �o�o�oO�o�o�o #5�oYk}�� �B�����1� C��g�y��������� P����	��-�?�Ώ c�u���������ϟ^� ���)�;�M�ܟq� ��������˯�O�O� �O�_$o6�H�m�l�~� ������"��������  �2�D�V�h�6oh��� ���������b�/�A� S�e�w߉�߭߿��� �������=�O�a� s���&�������� ����9�K�]�o��� ����4��������� #��GYk}�� 0����1 �U��ڿxϝ�� ����/ֿ(/&/ P/b/t/�/�/�/�/�/ ��??)?;?M?_?� �?�?�?�?�?�?l?O O%O7OIO[OmO�?�O �O�O�O�O�OzO_!_ 3_E_W_i_�O�_�_�_ �_�_�_�_�_o/oAo Soeowoo�o�o�o�o �o�o�o+=Oa s�@��v�/�/ ���&�8�J�\��� �z�����ȏڏ�� �"��/Y�k�}����� ��
ן�����1� C�ҟg�y��������� P����	��-�?�ί c�u���������Ͽ^� ���)�;�M�ܿq� �ϕϧϹ���Z���� �%�7�I�[���ߑ���ߵ����ߓw�t*default���=�*level�8��/�A�S��� �tpst[1]�U��y��tpi�o[23��t��u���4�Z����	menu7.gif�M
.�133�@�5H�h-�[�+�4o�u63� L�����������f� 3EWi{���������prim=.�page,74,1"@Yk}���6�class,13 ��� //$/��5*/`/r/�/�/�/��N/�/�/??*?-?18Fg?y?�?�?�?�/�6�?�?�?�O!O3O��$UI�_USERVIE�W 1�q�q�R 
�A�:O�mOO�m�O �O�O�O�O_�O3_E_ W_i_{__�_�_�_�_ �_�O�_oo�_Soeo wo�o�o>o�o�o�o�o �o=Oas� 0o���(��� '�9��]�o������� H�ɏۏ�����Ə 0�B���f�������ş ןz�����1�C�� g�y�������Z���ί �R��-�?�Q�c�� ��������Ͽῄ�� �)�;�M���Z�l�~� ��������ߤ�%� 7�I�[�m�ߑߣߵ� ���߄ώ���
�|�.� W�i�{���B����� �������/�A�S�e� w�"����������� +��Oas� ��L��� ��"4F���� ��l��/#/5/ �Y/k/}/�/�/LV/ �/�/D/�/?1?C?U? g?
?�?�?�?�?�?v? �?	OO-O?O�8