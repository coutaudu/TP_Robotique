��   ��A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_  �$$C�LASS  ������D��D�VIRTUAL�-9LOOR ���D?8�?���m8��M,  1 <dYH82 }~}���D'������ <i<?/Q/c/5/�/�/�-_ �/�/�/�+_�$MNU>A2">�� 	 8i	/ ��+?e?O?a?�?�? �?�?�?�?�?OO%O OO9O[O�OoO�O�O�O��O�O�	5NUM � ��>�>Pda�t2TOOL?�4 
';/u_DR �O�_�_�O�_�_�_�_ oo%oOo9o[o�ooo �o�o�o�o�o�o�o 9#EoXKQ+V[=9Vx.
