��   to�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����UI_CONF�IG_T  �$ 5$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY5]0�ODE�
1CWFOCA �2C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� �4 TOUCH�P{ROOMMO#{?$4 ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"��%�!BA�!j ?��"BG�%$PM��X_PKT�"I�HELP� MERޱBLNK$=EN�AB�!? SIPMoANUA� &�USTOM0 �t $} RT_OSPID�p4Cx4n*PAG� ?^�DEVICE�9S�CREuEF����7N�@$FLAG�@�
&�1 � h 	$PWD_ACCES� E �8�C�!~�%)$LABE� O	$Tz j�0�q!@D�	 [2US�RVI 1  < `� vB�nwAPRI�m� �U1�@TRIP�"m��$$CLA�0 �����A��Rz��R�@VIRTT1�O�@'2 )�7�)�@�R�	 �,��?���R�PSSQ�� ,/ �Y03_��
 ���Aw_�_�_�_�_�_�_ s_oo ,o>oPobo�_�o�o�o �o�o�ooo(: L^p�o���� ��}�$�6�H�Z� l��������Ə؏� ���� �2�D�V�h�z� 	�����ԟ����� �.�@�R�d�v���PTPTX�������� s �Ǖ���$/so�ftpart/g�enlink?h�elp=/md/�tpmenu.d�g��$�6�H�Z��&��pwd����� ˿ݿ���%�7�I� [��ϑϣϵ����� h�z��!�3�E�W�i�*?T��AMV/VS��($�ϻ������������AQ,�._��8����ߜ�lS�ْNQ��P���  a����Z@����f����*��Ca2 1��EPR \� }Y0REG VED������wholemo�d.htm"�si�ngl3�dou�bJ�trip�b�brows {�f������������ /Aj������/�dev.s8�lh�]�� 1�	t� ���e�5GY#�}������ �@//*/</N/`/`r/�/�/�/�& @/ �/�/�/??1? 6�� ��e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�Ow�O�O �O�O__1_C_U_g_ y_�_�_�_�_�_�_�_ 	oo-o�hozo�o�o �o�o�o�o�o
?. @!v�??Q?7o ������%�7� `�[�m��������Ǐ ������O��E�W� i�{�������ß՟� ����/�A�S�e�w� ��Woį֯����� 0�B�T�f�a����k� }�ҿ俛���,�'� 9�K�t�oρϓϼϷ� ��������#�L�G� Y�'�y�sߡ߳����� ������1�C�U�g� y���������ﳯ  �2�D�V�h�z����� ��������������. @��	������ ����%7 `[m����� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?�|?�? �?�?�?�?�?�?OO BOTO#O5O�O�O�J��$UI_TOP�MENU 1�u@�AR �
X�AT1)*default_?�H=	*leve�l0 *P ��O�5_4_F_�tpio[23]�tpst[1yX oP�O�_Z_S_�_�_��_�	menu5�.gif�
*a1I3/i(c1/k)b4/ko�Q��{o�o�o�o �o�o�oS2�o%7I [m���� ���!�3�E�W�i��{����prim�=*aclass,5��ÏՏ�������13�H�Z�l��~������page,153,1��@Ο��������8��O�a�s���������ͯ߯���L9 �@�A�OM�]?��Q=�wo��Vty�]r_�QOmf[0�_�\	���c[164yW�5�9yX�Qeo��A�#h2 Wo-m��CjOo9gVj�� �d-�?���0�B�T� ��xߊߜ߮�����a� ����,�>�P��ߡ�2b��������n� ���'�9�K�]����� 6���������������1��$6HZl�����ainedi�E������zwintp���(: L^pO6�A8�z� �V�_H����// ,/>/P/�_p/n/�/�/ �/�/�/�/?)?�oM? _?q?�?�?�?���?�? �?OO%O�?IO[OmO O�O�O�ODO�O�O�O _!_3_�OW_i_{_�_ �_�_@_�_�_�_oo /oAo�_eowo�o�o�o �oNo�o�o+= �oas�������5��Y�k���u�#?5�Ӻs��R�w�ſ_�u��*�,φ����@�Æ��.�|�R�6_�u7�����Ϸ�ɟ۟ ���V#�5�G�Y�k� }������ůׯ��������1	�G�Y� k�}�������ſ׿� ��Ϝ�1�C�U�g�y� �ϝ����������	�ߪϼ�6"�W�i�{�0�ߟ�����74���� �����#�G�Y� �/@����������� ��z��B�T�f�x� ��������6?��	 -?Q�u��� ���p); M_������ �l//%/7/I/[/ m/��/�/�/�/�/�/ z/?!?3?E?W?i?�/ �?�?�?�?�?�?�?�? O/OAOSOeOwO2�D� �Oh�2����O�O__ =_<_N_`_�Ol_�_�_ �_�_�_�_oo��Ko ]ooo�o�o�o�oO�o �o�o#5�oYk }���B��� ��1�C��g�y��� ������P����	�� -�?�Ώc�u������� ��ϟ^����)�;� M�ܟq���������˯ �O�O��O�_$o6�H� m�l�~�������"��� ����� �2�D�V�h� 6oh������������ b�/�A�S�e�w߉�� �߿���������� =�O�a�s���&�� ����������9�K� ]�o�������4����� ����#��GYk }��0���� 1�U��ڿx� �������/ ֿ(/&/P/b/t/�/�/ �/�/�/��??)?;? M?_?��?�?�?�?�? �?l?OO%O7OIO[O mO�?�O�O�O�O�O�O zO_!_3_E_W_i_�O �_�_�_�_�_�_�_�_ o/oAoSoeowoo�o �o�o�o�o�o�o+ =Oas�@�� v�/�/���&�8� J�\����z�����ȏ ڏ���"��/Y�k� }�������
ן��� ��1�C�ҟg�y��� ������P����	�� -�?�ίc�u������� ��Ͽ^����)�;� M�ܿqσϕϧϹ��� Z�����%�7�I�[� ��ߑߣߵ����ߓw��t*defau�lt��=�*level8��/�A�S���� tpst�[1]U��y��tpio[23��t��u��4�Z�����	menu7.gkif�
.�133�B@�5H�-�[�+�4o�u63�L��������� ��f�3EWi{ ��������prim=�.�page,74,1"Yk}����6class,13��� //$/��5*/`/r/�/�/�/��N/�/�/`??*?-?18F�g?y?�?�?�?�/�6��?�?�?O!O3O���$UI_USERVIEW 1�q��qR 
��:O�mOO�m�O�O�O�O�O_ �O3_E_W_i_{__�_ �_�_�_�_�O�_oo �_Soeowo�o�o>o�o �o�o�o�o=O as�0o���( ���'�9��]�o� ������H�ɏۏ��� ��Ə0�B���f��� ����şןz����� 1�C��g�y������� Z���ί�R��-�?� Q�c����������Ͽ ῄ���)�;�M��� Z�l�~��������� ߤ�%�7�I�[�m�� �ߣߵ����߄ώ��� 
�|�.�W�i�{��� B������������/� A�S�e�w�"������ �����+��O as���L�� ���"4F� �����l�� /#/5/�Y/k/}/�/ �/LV/�/�/D/�/? 1?C?U?g?
?�?�?�? �?�?v?�?	OO-O?O �8