��   to�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����UI_CONF�IG_T  �$ 5$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY5]0�ODE�
1CWFOCA �2C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� �4 TOUCH�P{ROOMMO#{?$4 ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"��%�!BA�!j ?��"BG�%$PM��X_PKT�"I�HELP� MERޱBLNK$=EN�AB�!? SIPMoANUA� &�USTOM0 �t $} RT_OSPID�p4Cx4n*PAG� ?^�DEVICE�9S�CREuEF����7N�@$FLA�G�@[2�1 � h 	$PWD?_ACCES� E �8�C�!�%�)$LABE� '	$Tz j�0q!�@D�	 [2USR�VI 1  < 	`� vB�wA7PRI�m� U1ޖ@TRIP�"m��$$CLA�0 O����A��R��=R�@VIRTT1�O��@'2 )�7)��@�R�	 ,R��?���RP�SSQ�� , ��Y03_��
 ���Aw_�_�_�_�_�_�_ s_oo,o >oPobo�_�o�o�o�o �o�ooo(:L ^p�o����� �}�$�6�H�Z�l� �������Ə؏��� �� �2�D�V�h�z�	� ����ԟ�������.�@�R�d�v���P?TPTX�������� s ������$/sof�tpart/ge�nlink?he�lp=/md/t�pmenu.dg@��$�6�H�Z��&��pwd�����˿ ݿ���%�7�I�[� �ϑϣϵ�����h� z��!�3�E�W�i�?T��AMV/VS��($�ϻ������������AQ,�._��8����ߜ�lS��NQ���P���  �����Z@����f�p��*��Ca2 1�E~PR \ �}Y0RE�G VED������wholemod�.htm"�sin�gl3�doub~J�tripb�brows{� f������������ /Aj�����/�_dev.s8�l�4]�� 1�	t��� �e�5GY#}�������  �@//*/</N/`/r/0�/�/�/�& @/�/ �/�/??1? 6��� �e?w?�?�?�?�?�? �?�?OO+O=OOOaO sO�O�O�Ow�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_	o o-o�hozo�o�o�o �o�o�o�o
?.@ !v�??Q?7o� �����%�7�`� [�m��������Ǐ�� ����O��E�W�i� {�������ß՟��� ��/�A�S�e�w��� Woį֯�����0� B�T�f�a����k�}� ҿ俛���,�'�9� K�t�oρϓϼϷ��� ������#�L�G�Y� '�y�sߡ߳������� ����1�C�U�g�y� ���������ﳯ � 2�D�V�h�z������� ������������.@ ��	������� ���%7` [m������ ��/!/3/E/W/i/ {/�/�/�/�/�/�/�/ ??/?A?�|?�?�? �?�?�?�?�?OO�BOTO#O5O�O�O�J��$UI_TOPMENU 1u@��AR 
�X�AT1)*d?efault_?H=�	*levelw0 *P �O��5_4_F_�tp�io[23]�?tpst[1yXoP �O�_Z_S_�_�_�_��	menu5.�gif�
*a13$/i(c1/k)b4/ko�Q��{o�o�o�o�o �o�oS2�o%7I[ m����� ��!�3�E�W�i�{�����prim=�*aclass,5���ÏՏ�������13�H�Z�l�~�������page?,153,1��Ο���������8 ��O�a�s��������@ͯ߯���L9�@ �A�OM�]?��Q=�wo���Vty�]r_�Qm�f[0�_�\	��c�[164yW�59@yX�Qeo��A�#h2Wo -m��CjOo9gVj�ϊd -�?���0�B�T߫� xߊߜ߮�����a��߀��,�>�P��ߡ�2 b��������n﬏ �'�9�K�]�����6����������������1���$6HZl��~��ainediE�������zwintp���(:L ^pO6�A8�z��V �_H����//,/ >/P/�_p/n/�/�/�/ �/�/�/?)?�oM?_? q?�?�?�?���?�?�? OO%O�?IO[OmOO �O�O�ODO�O�O�O_ !_3_�OW_i_{_�_�_ �_@_�_�_�_oo/o Ao�_eowo�o�o�o�o No�o�o+=�o as�������5��Y�k���u�#?5�Ӻs��R�w�ſ_�u��*�,φ�����à���.�|�R�6_�u7�����Ϸ�ɟ۟� ��V#�5�G�Y�k�}� �����ůׯ����
����1	�G�Y�k� }�������ſ׿��� Ϝ�1�C�U�g�yϋ� �����������	���ϼ�6"�W�i�{ߍ�������74������ ���#�G�Y��/ @������������ �z��B�T�f�x��� ������6?��	- ?Q�u���� ��p);M _������� l//%/7/I/[/m/ ��/�/�/�/�/�/z/ ?!?3?E?W?i?�/�? �?�?�?�?�?�?�?O /OAOSOeOwO2�D�O h�2����O�O__=_ <_N_`_�Ol_�_�_�_ �_�_�_oo��Ko]o oo�o�o�o�oO�o�o �o#5�oYk} ���B���� �1�C��g�y����� ����P����	��-� ?�Ώc�u��������� ϟ^����)�;�M� ܟq���������˯�O �O��O�_$o6�H�m� l�~�������"����� ��� �2�D�V�h�6o h������������b� /�A�S�e�w߉�߭� �����������=� O�a�s���&���� ��������9�K�]� o�������4������� ��#��GYk} ��0���� 1�U��ڿxϝ ������/ֿ (/&/P/b/t/�/�/�/ �/�/��??)?;?M? _?��?�?�?�?�?�? l?OO%O7OIO[OmO �?�O�O�O�O�O�OzO _!_3_E_W_i_�O�_ �_�_�_�_�_�_�_o /oAoSoeowoo�o�o �o�o�o�o�o+= Oas�@��v �/�/���&�8�J� \����z�����ȏڏ ���"��/Y�k�}� ������
ן���� �1�C�ҟg�y����� ����P����	��-� ?�ίc�u��������� Ͽ^����)�;�M� ܿqσϕϧϹ���Z� ����%�7�I�[��� ߑߣߵ����ߓw�t�*defaul�t��=�*level8��/�A�S���� tpst[�1]U��y��t?pio[23��t�u��4�Z����	�menu7.gi5f�
.�133�@��5H�-�[�+�4o�u63�L����������� f�3EWi{� �����~�prim=.��page,74,1"Yk}����6class,13��� //$/��5*/`/r/�/�/�/��N/�/�/?0?*?-?18Fg?@y?�?�?�?�/�6�?��?�?O!O3O��$�UI_USERV?IEW 1�q�q�R 
��:O�mOO�m�O�O�O�O�O_�O 3_E_W_i_{__�_�_ �_�_�_�O�_oo�_ Soeowo�o�o>o�o�o �o�o�o=Oa s�0o���(� ��'�9��]�o��� ����H�ɏۏ���� �Ə0�B���f����� ��şןz�����1� C��g�y�������Z� ��ί�R��-�?�Q� c����������Ͽ� ����)�;�M���Z� l�~���������� ��%�7�I�[�m�ߑ� �ߵ����߄ώ���
� |�.�W�i�{���B� �����������/�A� S�e�w�"������� ����+��Oa s���L��� ��"4F�� ����l��/ #/5/�Y/k/}/�/�/ LV/�/�/D/�/?1? C?U?g?
?�?�?�?�? �?v?�?	OO-O?O�8