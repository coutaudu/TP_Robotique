��   ��A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ��	��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !� FTP�_CTRL. =@� LOG_8	��CMO>$DN�LD_FILTE�R�SUBDIR�CAP���HOv��NT. 4� �H�9ADDRT�YP� A H� NGcTHOG��z �+LS/ D �$ROBOTI<G BPEER�� �MASK@MRUv~OMGDEVK���RCM+ � $�x� ��QSIZN�TIM$ST�ATUS_�?MAILSERV��LANT� =$L�IN�=$CLU���f=$TOcQ�$CC5&FR5&A�LAR�B�TP��\#VARd(�R�DM*� $D�IS� �T�CPIo/ 3 �$ARP�)_IPFOW_��oF_INFA~�LASS�HO�_� INFOz"T;ELs P~����� WORD�  $ACC�E� LV��OU| wORT ��ICEUS 0 �  �$�#  ����r1��
���
g0VIRTU�ALo?�1'0 �5/
���F��d02���4�5���� �=��!y1O����$ETH_FLT�R  �6�3 *��������K��� �=2K�"SHA�R� 1�9 # P O�O�4�O�O �O_�O*_�ON__Z_ 5_�_�_k_�_�_�_�_ o�_8o�_ono1o�o Uo�oyo�o�o�o�o 4�oX|?u� �������*� �S�x�;���_����� 䏧��ˏݏ>��b� %���I���m������ �ǟ(��L��E����q���i�ʯGz _L�IST 11Mx/!1.�0ӯ����1���2551.M������5�2
����0�B�T�f�x�3���������̿޿x�4���q� �2�D�V�x�5r�������ϼ���x�6���a� �"�4�F� ���1��K��}0� 'Q����=��1� C��g�y��^������Q��������9� K�]�o�.���������0J$� �>�$�%� ��=� �6�5	1�:�9�@@H!� X���rj3_t�pd���1 �0y1!KC�0�m	��<�6�!CP0�����!CO�Nn03nzsmon�