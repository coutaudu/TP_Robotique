��   ��A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ��	��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !� FTP�_CTRL. =@� LOG_8	��CMO>$DN�LD_FILTE�R�SUBDIR�CAP� HOv��NT. 4� �H�9ADDRT�YP� A H� NG#THOG��z +�LS/ D $ROBOTIG �BPEER�� MwASK@MRU~;OMGDEVK%�RCM+ �� $�� ��QwSIZNTIM�$STATUS�_�?MAILS�ERV�LANT�� =$LIN�=�$CLU��f=${TOcQ$CC5&{FR5&ALAR��B�TP�\#VA�Rd(�RDM*>� $DIS�%OTCPIo/ 3 �$ARP�)_7IPFOW_�޳F_INFA�~LASS�H{O_� INFOz"wTELs P~���� WOR�D  $AC�CE� LV��O�U wORT >�ICEUS 0���$�#  �S��r1��
��
g0VIRTUALo?��1'0 �5
���F����%�2�5��� �=���!y1O���$ET�H_FLTR  \�6�3 ���������K�� �=2�K�"SHAR� 1}�9  P O�O�4�O�O�O_�O *_�ON__Z_5_�_�_ k_�_�_�_�_o�_8o �_ono1o�oUo�oyo �o�o�o�o4�oX |?u���� ����*��S�x� ;���_�����䏧�� ˏݏ>��b�%���I� ��m�������ǟ(� �L��E���q���i��ʯGz _LIST� 11Mx!1E.�0ӯ���1�>��255.M��&����5�2
��@��0�B�T�f�x�3����������̿޿x�4 ���q� �2�D�V�x�5r�����Ϫϼ���x�6���a��"�4�dF� ���1�K���}0� Q����=��1�C��g�@y��^������Q�� ������9�K�]�o� .���������J$� �>�$�%� �=� �6P�5	1��9�@@�H!� X��rj3_tpd����1 �0y1!K�C�0�m	���6�!CP0����?!CONn03znzsmon�