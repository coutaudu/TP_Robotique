��  �\�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A9  �����ABSPOS_�GRP_T  �  $PAR�AM  ����ALRM_R�ECOV1  � $ALMOEkNB��]ONi�I M_IF1 �D $ENAB�LE k LAS{T_^  d�uU�K}MAX� �$LDEBUG�@  
0���APCOUPLE�D1 $[PP�_PROCES0S � �1�G�PCUREQ1� � $SOF�T; T_ID�TOTAL_EQ� �$,NO/P�S_SPI_IN[DE��$DX��SCREEN_NAME �/SIGNj���&PK_FI� 	$THKY��PANE7  �	$DUMMY1U2� �3�4�~GRG_STR1� � $TI�T�$I��1�&�$�$�$5�&6&7&8&9'0''�%!'�T%5'1?'1I'1S'�1]'2h"GSBN�_CFG1  �8 $CNV_�JNT_* �DATA_CMNT�!$FLAGSL�*CHECK���AT_CELLS�ETUP  �P� HOME_I�O� %:3MA�CROF2REPR�O8�DRUNCD̻i2SMp5H UT�OBACKU0� �	DEV�IC#TIh�k$DFD�ST��0B 3$INTE�RVAL�DIS?P_UNIT��0w_DO�6ERR�9�FR_Fa�IN^GRES�!Y0�Q_�3t4C_WAx�4�12JOFF_� �N�3DEL_HLO�G�2�jA�2?�1k@�?�� ��ՁH X_D�#	� d $CARD_EXIST��$FSSB_T�YPi� CHKBoD_SE�5AGN �G� $SL?OT_NUMZ�AOPREVD�G ��1_EDIT1
� � h1G=�H0S?@f%$EP<Y$OPc �iAETE_OK��BUS�P_CR��A$�4JVAZ0LACIwY1�R�@|k �1COMMEc@$D�V�QO�k@:Y��$QL*O�U/R , $��1V1AB0~ O�L#eR"2CF�D X $GR� z� S!1$MB_@NFLIC�3\`
�UIREs3��AO}MqWITCHWc/AX_N.0S�=`�_;G0 � 
$WARNM'@0f��@� LI? �a�NST� CORN���1FLTR�eT�RAT@0T�` �0ACC�1�` |�rORI�P�Cxk;RTq0_SF� �!�CHGI1 E[ TT`u3I*p�TY�2QqK*2  x �`� 1�B.*HDR�J* ���q2�v3�v4�v5��v6�v7�v8�v9�#QCO�$ <�� Mo_oqh�s1<`O�_MOR. �t 0Ev�N5G� �0BA� �Q�t�Q}��r��@��v���P�0����h�`^P/P�2н �p�Jp_R�bLq�@�J	r	�$�JV�@�CD��m|g�v�uMtP_}0OFܚ �  @� RO1_����aIT8C��ONOM_�0�1��pq3W ���$ �����|hP���mEX �`G�0� �0"��`�b�
$TFR�J �DM3��TO�3&@U=0^�� ��H�2��T1m�E��� ��e��f��f��0C�PDBGDE�m�@$`PU�3�f)����AX 1�dbETAI�3BUF�F�����!� � ˧�`P�I���PL�M�K�MX���[�FL�S�IMQS��KEE��PAT�`�!�� �����MCU�5 �$}1JB�`-��}1DEC㺋��܂�S� �7PCH�NS_EMPvr#$GA�'��@_y�q3��`1_FP͔x�TCR�SPEubw�q0 �cg�S�!�� V�A����!����JR!0��SEGFRApv r�}R�T_LIN�C��PVF�������Y��P��)B|��وD )\� }f�e	�"��	��.0��Z��Ql��SI!ZCuх�d�To�A���ڭ�	�RSINF ��p����?���ܭ���s���LItx�1��gCRC�eFCCC�`���>�R��mRM�Al�R��P� �$�DȆd�c��C��j@TA������@��l���EVT���jF��_��Fw�N�� ��f��!�� B2���������1C���! ����hRG�Ps�
qF��7bg�qD���2g�LEW(��s� �e�>�P�|+�C� ��&�pou2|��A6NHwANCI�$LG�`�-��1�Pd��@�d�aA?@l���~0R��z�j�ME��uAk��eRAs3jAZC���:T�OEqFCT�q����`F�`m�g�̰�ADI;� q�� �l��`��`�`|�H�S0=P�r��AMP�Ĥ��Y8C?�MAESЈ���r�I�$�  *�I���GCSX�a�!�p�	$JTpT�X�C�_ N�@h�IMG_�HEIGH�A�W3ID��h�VTE��U�0F_A��- ��@EXP(�c-%��CU���QU�1 �$`TIT�1�9RISG1ꀿ��DBOPXWO���0 zp�$SK���2ԑD�BT% TR�@ 	!^�Q0TC�� `���DJ�4LAY_C�AL�1iR� '�'P1L	3&@�0ED���'�Q�'�Q�Py ��!�"�"1�PR� �
� �q��!# lT A$wq$��
�L@9$M?_3Gp� )%s?�4C�!&�?�4gENE�ax�'�?�_3!0RE�`�2(�H C�p #$LC$$@3�B� hK��VOa _D6G�ROS�bcvh�D���AMCRIGGER�eFPAyS���ET�URNcBo�MR_�o�TU�`)�2@EkWM����GN`���CBLA���EΑ<�P��&$P� 9�#'�@�QU�C�D���0DO����-DAS��3FGO_AWAYFCBMO���Qm� �CSC0EVI>@ �) HJ`1vRB�w���SPIhpJ�SyP`wVI_BY��|S�UHSL�r*XP�$��avVTOFB�\�dFE=A1v�SvT�HS�+ 8��D1O?��cnpMC%�d��P��)b�R�& `�,� $���J  �c #fc ��faסߠebit�cH�fa�"af9Wr��dNTV�fbV-pr���؃���g�s�?�J�?��0��SAsFE̕v_SVq��EXCLU�!��N��ONL+�<sY�T�ktOT!!��HI_�V5�PPLY_`,�etw�]fjs_M8�� $VRFY	_�#�O�� �v!�1��s�bFc"�Q #-�0� ~�_�:�� CeSG� .�
$���@�A�����U�REV0�-�$��UN�0x K�vU��턍��@���l�i�!q����"EF�f`I�2/��$F�N�X$�OT�@jS?$DUMMY
1ׄ�1ׄ����M�PNIG20 L����4�r��A`a�DAY҆e`ADiT� ��؃5F��EF $���1�0�ѧ�Y�_3� _RwTRQݑ2 D_�-Ot@RQ:���'�<��Y� 21�����~�jT|��s�¡3 0��ؑ�	�גS��U�@��"CAB�¡4����$��$ID��PW��ӕH�g�ViWV_Ӑ��0��DIAG�q¡5?� $$V�@a�T�ǃ���� ��
0	�R�25��VE� J�SW������(����~���2ZP~�OH̔��PP���IRs!	�B��7�����A8ᇀ��BAS9q�@z ���iV���4���Cנ�RQDW&�MS9���A����<���LIFE� ����10��N��
�ɵ@i���
���^Ui�Cm+7QN�@Y����gFLATj�OV6�նHE���UPPIO��w��� _6�p� , �6 `�pCACHE-�m���Es�B�SUFFIX�e`� ��@��R�؃6���!MSW��7bKEYIMAG�CTM%AH���<�A��INPURę �OCVIEʠ�!8 h�� L�d��c�?� 	�!"�9~��$HOST� !R�
0Z�0Z�G��Z�R�Z�EMAILp\ E�� SBL���ULG2:"҃�C�OU��T�T�0y�;� $��eS�Ӑ4�IT1cBUF@ǂa�NTf j 5�	B��mTC�dA��s#���SAV<��҅�E@K@b2W�Ppm�PC�e�0ˤ��_��"�`F��OTRBu�?P�p�M�e���r��Z͓D�YN_�� <��DHtU� �U���_TR_IFS�W�8O��A�!=0��/�p�Ӡ�#$@TIKYD#&�L�A����K����/�DSP��/�PC��IM<���sM�w�Uf�+�XE�p��I�P�c/���D0��T!H0�|�TLA���HS��ABSC$H���F��s�dk�$���oSCi�ʖ�1�!ڤ!>bFUI�DU���c��@PE���C�D�	 ���W�R_�NOAUTO�!?���$���:�PUS�C0�C�"�s��!��� @H *�LI ��� jUs@�c>
1< 1<G�<R�<��<798999��;�E1R1_1l1�y1�1�1�1�2���GR`�H�l2y2�2�2��2�3�3E3TR_3l3y3�U3�3�3�4��XTz�NaA <���� �]V �jU�7���FDRi�BT ��	���pò�17òREM��9FQ̲OVMb��5�A�9TROV�9D�TG�JMX#LINp�98PJf�IND2@�ʲ
^H* s�$DG
�X+�@M`ɵ��9D��@RIV�U̲oGEARb�IO��	K�2ʴN$��HY����_p�`�a̲Z_MCaM��ñ�0,�URw�C ,�Wq?�  �p?0P��K?0QEop8Q�1&�`COԐO`D��n�5P1av�RI�QTnz�UP2�pE G���TD��os�S0�HQp�W�Ud1��BAC��F TP����Ł)
]qG�U%��� t IFI�� XP]`+���UPT̢CaFMRE2�5G���1�s�2LIxaFc�7�O�O�OPF��ʵ�2_��N"��_�����M�F�O��MDGCLF�D7GDYxLDHQ�DA5Ѷ�Oɴ'cE�Hl ��i T�FS��F�I P��xqL`|
�s�$EX_wq��xwq1��EZwq3z�{5�v�GRA�Pθ4J ��tSW�%�Ot�DEBUG��#���GR0���UnZBKUe O1 7 PPO`0�b�CԐ�t�MS�`�OO��^�SM�`E�K⦁��0_E �K S��Pv��T�ERM��L��Ҁ�'ORI`��M�����SM_�P�҅�N\�����TAǉO����UP�P� 9- ��2K$����L$SEG�%pE�LTO��$US]ED�NFI�<��Pt�� ��
�M$UFR�R��� 6����&�`OT��pT���0NST��PATxx���PTHJI� EH�s� �=�AR���I���V��<�REyL�r�SHFT �=���ۘ_SH:�M�O�Ɔ р��5�O�a�0OVR��r�&��I��dU� ^�AQY��Q`��ID�MhSp�� q� ERVD x�7 &�h2������!0`ӥ�!`RCXQrŏASYM"�r�=�WJP�h1d@EhSב�����U'�������ф��P����V�OeR��M@c��GRo��tQ���U���l����W�S�E�R � �h�QTOC6�:�Q��OPbm���(*tv��1OA�KRE��RT�r�O
�,]⮒e�R��>�����Te$PWRf�@IM0ũ�R_���S�]� S�P�$H�U[�_ADDR�6Hr�G�������vѷR=p��8�T H�pS` ���#���#0��_��lSEkq���S� �sU $���_Dm0=���+һPR����T�T��UTH7�V }(� OBJECa�!(Q�Q$�6LER��_�8�W�px7���AB__A�Գ�S|��I�DBGLV��wKRLp�HITE�[BGD�LO����TEM���%B�g��SS�@7�HW��C���X��\�I�NCPU�rVISIOR���Di���j���j�l �IOLUN��Y} �@C��$SL��$I�NPUT_u�$�0���P�@���SL�p��Z������I�O@�F_AS]r[�P$L�P���Q-�".Uƀ)�T��� ���z�HY�7T�-�d1��UOPZu\ ` �r�6BBD�B@K���B�P90�����K�����d1UJ�6] �� �PNEV�JO�Gk���DISBcJ�7/�OF�$J8�	7W IT�'97_LAB���) Q�APHI�`Qt(mDypJ7J���0�p_KEY�`� �Kk��0\s^� �@��V��{6�C�TR퓵FLAG��rLGʴ_ ��9`y8���sLG_SIZ�ԧPXp�FDI"Q� 
��	�� Xp���9����2@SCH_H��R�R� N�r`~���@�p�q��1�`UH�����L#�DAU%EAP�k�ܴ3") �GHݲ�OGB�OO�Rat B3��IT�3g$�`/��REC|*SCRN,� /�DI.�Sl�=pRGMb�0�,��'���H�"���S���W�$��$'�JGM7MgNCHF�'�FN��6K;7PRG99UqFG8W�G8FWDG8�HL~9STPG:V`G8`G8n G8RS�9Ho�c;$�CY��3&�'��p�'IUG�[4�' H��&� <�N2G+9�PPORG�:�%�3P/6�OC$�J8EX#�TKUI95Ii�#�B �#�C3�C70;11���`AC�'1��!NO�F�ANA�6��`VA�IQ ��CL�a��DCS_HI	�NR��bMROSX�aVTSIxWrjXSvX�(IGN"���481�  `UUDE�V$��BU`��bj� _�T�B$#EM�[��T �
��c� _���e�W�TQ`m@19e29e39aq@�T}Q��d ������{�5���%��ID opX�.�4�=a�&���f+STs�R4 Y�p1�~�` c$E�fC�k�Б��f�f���D��e LL�B��pW� )�� �C����PЄ���"�#_ f �:��V����!�s|�C��g ���CL�DPs���TRQL�Ii � �y�tFLAG�b�p�a�s=QD���w=�LD�u�t�uORG �2�r���8���ç�ҙt0�h �C 	�u�5�t�uS���T�p� s�!���>��RCLMC��<�`N���������MI�Ν�i d�yaRQz� s�DSTB��Ɯ` ��!'�AX���� *�C�EXCE�S���MO���j�P�������Nџ�5k���_A���Я�A�S��pKʴl q\L��$MB>��LIw��REQU�IRˢ
��O�D�EBU`B��LSpM�m��4�Z���������ND	!ǰ��n0�����DC�B$INeЫ!$�� ��¢PN�b�C�PS�T�� o��LO�C|fRI&�|eEX��A��}a���OD�AQ�p
�$ON�RMF�@`���iRrJ@\u����SkUP����FX��IGGz! q �s�Rs���RsFRtR��%�cιs�޸�s��ΐ<�DATAg*�Eq�E��T��N�Rr tN�MD
K�Ix�)YƎPd��a�H/�"dĸ�Ue�ANSW�!d�a�A
d�D&�);��󔀟зs ��CU"V����p7�RR2��t����Z���A�� d$CALI �ҝGAQ
�2��RI�NP0�<$R�S�W0ʄH�y�ABC~_�D_J2SE4�\�X�_J3s�
m�G1SP?�< �Pm�B��3���������qJy��Մ�V_O�Q�IMy���CSKP �z��:S�J<!���Q�3��3�)�$�_cAZ����e�EL�Q�����INTE��"bu����7���%p_N��v����ah���䛒w��DI{�F��DHc�����x� �$Vв��a$;1$ZbN`b������yH ��$S v�TqACCEL�QU�ׁd�WIRC��T?�yT�a�c$PSc��rL  & ���s���z��BP{�PATHZ���p���3���f��_6a$� ��M`Cܴ�k�_MG�!$�DD${�"$FW��=�`�@p�k�5�DE^PPABN���ROTSPEE�:a��p)�:aDE�F!�k��$USSE_�SP��CO@�SY� 6� ��YN �A� ���{��7MOU!NGO� sOL��INC�Ā,�]D'�=��(�ENCS�#����k�,%���IN�bI��>���)�VE"Ӡ�23_U�b�LOWL�QI@���pi�D,@�����Wp�i��C���MOS��PӔMOܰ����P�ERCH  �OV� �1'|a<#�a� ���a2�m"�,����$P��A��%LT�ӀЗ�ך����&�T�RKE$�bAYLOA���"�� 1��538-��`S�RTI��K�`MOM�B'���2����\
�3��9b�5�DU����S_BCKLSH_C�� �5&D ��°4dx�:+�CLAL`����A0���5CHKt�p�eSRTY�@@(��@�e$�<�_�cN$_UM��=ICJC�$SCLWD� LMT��_L6���pE��|GEvM�@�Ku@���E����Ц1
� �Du(P	CB!u(HYp;�(@E�C��]rXTk�6C�N_%�N�S7V׃S�P� g(V��c|V�Q��{UXC!`HMSH�c%�6l$�{1{��2���U��$PALGD;_PFE*3_�p�d@6% �q3)dEJaGxpy�c�OG*W>n2TORQU� �� # 9l ��"o1l �b_WY5 4_�e�e�eI�kI�kI�FE��a��x]�. �VCZ�0!��"r1�(~u�<2�/uJRK�(|mr`v��DBL_�SM7��M��_D9L�GRV�d�t0�t�qH_�S�s���zCOS�{/0�xLNop
�+u�������aH�6��a�uZ�&�qMY����r�TH�}��THET=0�NK23�тl��CBֆCB�C �h����d	��	��ֆSB�'��GT	S���C��,��S&���PS�6�`�E�$DU@И��
�G�������]1Q�2�$NE䗰I�(C�2R���	$��ŁAɅ����u�x�qLPH�uВ�ВS'�C�6�C�E�В�T�m�W�t���V�V�	��,�V;�VH�V�V�Vd�Vr�V��V��H�-�3�+��QJ��H�HV�Hd�Hr�H���H��O�O�OT��*�O;�OH�OV�UOd�Or�O��Ot��FВ��R�6�W��S�PBALANCEl���ALE>�H_ɅSP��'���6���E�PFULC���½����E���1uLUT�O_@=eT1T2�V�2N�1q�)�6Ԁ��:1�������U1T�� O{�c�`INSsEGq��REV���DIF�%��1�v����1w� OB���1�sg72x`)�A~�tLCHWAR���AB�Qi5$MECH�����(FAX1P�D,�����x 
-�aO�|7ROB% CR��o�z!R,��MSK_���9�z P !�_�� RV����$1 zR�����4�����IN|��MTC�OM_Cp=�{ �  ��v$ONORE��������| 4�`GR܌b�FLA|�$?XYZ_DA�B`^��DEBU?� ��$�} ��$�C;OD�1 o�>2��90$BUF/INDX� ����MOR��~ H ��W0e��6��5�4��J�&Q��@�TA���g2G��� � $SIMUL'`v�X#<�#OBJE���ADJUS1$ A�Y_I>az(DRO�UTG`>�W0_F-I=��T�`�	 ��I��Ф`� ���t���%D� FRI�3��T�5ROg`�E|�a� �OPWOnp���,|�SYS�BU⠙�$SOP����1U��PgRUN��<PA��!D;�s _m �B�1��ABc��@m I�MAG�1�ฐPf��IM��IN�p�d�RGOVRD�- oPq�xP��L_	ЄQ�<BWP�RBXP���AMC�_ED��� �@N��M"�A�0MY119�A��SL������ x $OV�SL[�SDI� D�EX@SR&OS�!p"V�`m%Nw!�aj� u#Њ'�(%"AQ0$_SsET�`��� @�`��"6�1RI�0
B�&_��'�!�!	�ฦ�/ lP ���T��<`ATUS~0$TRC��� ��/3'BTM87"1IY#$�4�A3 ��� DB��EmV",2�E���-1�� �0-1EXE�30)A!�2�2f4�#��� ��20UPI�19$�ИXNNX7qx#$q[9 �PG���� � $SU�B!16��!!1�#JM/PWAI�PPz#9E�LOy@9��$�RCVFAIL_C��RP<AR�  �)��QjPATs��E��R_{PL�#DBTB<a�nRRPBWD~F�UMl`�DIGT�<��[�ADEFSP>H� � L��3���@_�@7�CUNIr]7�@�1R�0�r�pk_L��P+1��	P����k�e`�qЭ J���N��KEQT@R�`W�HPP�B�� hB ARSIZE�P:� I�Q�S/ OR�#FORgMAT��DCO5 ,�Q~�EM%��T#S�UX� �"FQLI��B��  $>��P_SWI�д%�qp�@�@AL_ G� $�A���B!���C��DY$E6�1�,`C_�A� � �@�d���(aJ3r����TI�A4�i5�i6��MOM��c�c�c�c�c��BP@AD�c�f�cl�f�cPU
�NR�d�u�cu�b���R�� C$PIǖ oe��od�tWu�sWu�s Wu��vm{ �r�[!P��j!{�$�6�SPEED��Gb�tQE �D�v�DQE�@� �v���x�A��AQESAM�����Z��w[�QEMOV�򊔉��Л�����$���@1�䶄2���  ��`��%`�H<Т�IN�%`>������QB�2�	�2�R�GA�MM~Ʒ�I�$G#ET���;D_d��=
1�LIBR�1Gr]IT�$HI�0_�H;0��ǖE��ԘAΞ��LWɝ���p3��[b%�MTN+a�C�E����  ?$PDCK�$�;_=�� ��$bph$a�؅���c���f��)c _�$I� R"��D�����1rD��LE@����!�[h�n`MSWFLY��T�����Pq�UR_�SCR�3`�-�#S_SAVE_D�,~��3NO_`C�!�2 `d~���ojXv��qy ��0��ۻN���v� ̀Ja` <����љ��� �����x�v��|� x�6Û��1ERL����ߏ � ��YL Qs��؇Pу�ɣ�Ǟc����W������A�p�����M��(�CL'�(aC&"l�8"&�q/!PLMo���?� � $���g$W~���NG� ya~�8d|�?d|�Fd|� Md�@��᪐c�%`%X9POGc$aZ��P@ �� pB ��ʣUv��ҿ�����:_a_�� |B oi ~��i��c��c~��j����jE@ ���#��JU��\�z`��P�Q��PM� QU_� �� 8TPQCO�U̡^ QTH��H�O��c�HYS�PES��b�UEN�t��P}Od�   ��̽��"UN40*� �
@O���� P����oE`�}3GrRO�GRAG1��2�4O�����R���INFO�� ���� ����FQOI#� =(R�SLEQ�vK �uK �����D>@�������O�����s�ƑE�NU��A�UT���COPY����0�j!��M�N�� �m�C� �QR�GADJ�ᚓRX�R$9P.�.W,P,$�.�s�&CEX�@YC���FQRGNSD�� � $ALG�Oz���NYQ_FREQ��W=��v��T�#LA��ѫc=��uCRE�0�#� �IF�"��NAc�%�_G�&3(%���ELE-@ ��jbENAB�ҡPEASI_!|���N"@�q���&cBՀ��I �����qf�_`��"AIB�!K`E���pV��'BASUb�%����8�0���0$�!6�PUG$�� X� �" 2� ����>62=7;QX�ޠR5i6ER�-P�F��RGRIDd�13CB�P�wTY`#N�OTO�`��@���_$!Z�2C$O� ������[@P�ORqC�3Cv�2SReV )	DFDI�P�T_�p#@5D��?G3�=I"P?G5=I6=I7�=I8!A�F����~��$VALU�#�q�r$n��C��|C [%�����3!�n��PANp�vS0 R�0�Qn�TOeP`���$SPW�I�1:TR�EGEN8ZMROcX�7�s�v���FI�TR�#1B8Q_St��WMP��#Vѵq�U�q<!GRTb�Q�Slì� nSV_H�0DAY��P�PS_Y�����mSo�ARY�2�+0�CONFIG_SE_�PBn�d2���G�5� 4W�?�vv[δ6�PS~��� =@W�MC_Fl�|�a�L�~��SM����a�bNs����ܟc� ,R�FL��Г���YN�`|M�f0C���9PU��L�Y�ᦛ�DELA44pb�Y��ADY� �QSKIP�ŧ� ľ���O��N1T��o1^pP_���� }w`��ҵ��w�Q�y�Q �yV@�zc@�zp@�z}@��z�@�z�@�z9�q��J2Rf���fbEX��T�C�n�C���0rC���q�RD]C֩ ���R� ��M�ͅ����f�w�RGEA�R� ]��0E�D��ڝ�ER�a^�9C~UM_C�p�?J2TH2N��4�� 1� t�EuFI�1�� l(��4�\#����TPE���DO�]��� ��T���O3S���Ւ��(~��&�2.��4�F��X�j�|�����3.�����ß՟������4.��.�@�R�d�v���
��5.������ϯ�(����6.��(�:��L�^�p�����7.�������ɿۿ�����8.��"�4�F�X�j�|�^��SMSK��#��
�'�bPD�#�RESMO& ���f`瀘6�V4�IOT�I����B%�POWER�� 6�pa�����S ��e��$DSB� �!T/pyC�t�S232:���� *�DEVI�CEU�". t�RP�ARITY�.!OP�BITSFLOW0`TR�� R+P���R�CU��r UXT�ASK�RINx�F�AC��1"��� ��C�H���b�`_sC2����POM�tbPGET_�@�b� 8g0��1RSP[��߸� !��$USAp�1���� O�`� ��'`���_ON�P����'WRK����D�P�~��FRIEND 1x $UF��#w��TOOL~�MYH��`t�LENGTHw_VT��FIRM`ȧ��U E�е�UFwINV ��RGI�MAIT�I�r��Xzq�� G2 �G1�1U���d+�0_y�|O_�� ����#� ����@�TCs��D� �QG߀1#b`��`�� ���bo
�.%�S0#�R� �������XS ��v0L�T�H�0��&����)$IW�0�EDRpLOCK6'Aqwp�Q�Ui�Q$�20����4�.�:�1F�5�2*8�2�38�3F�� �G��!�����S��R�SV�P��VVV@(�`b`���b� �so:�|+e p�q	P]P�! ��S��U�d���A9@�'PR�P�&��SS�q� �q/����2� 0�0�20�haV#������E �U�{r
��S���� �c!RAQ{2�$P`N��`�BHA�n�L��rw2THI�C.� papC��T�FEREN1t5I�@H.�w1I8��3��K0G1�(�4���9�r���6_JFGP�R�`}q�b�C� �<q� *R }r�C 8�-F{� ��҆a�  2� �S�x����	d �$��Du��E�C$Pn4�CDSP�FJOG��P�p`_P�q:�O��1Fu��� L�KEPF��IR�A�D]`M&UAP&�E�%P��4�S`�@�R�PG:VBRK`�5�0:n0I��  aR�c�lR�Br A�R�C�@B�SOC�FJ�N�UD�#`Y15�q$S}VDE_OP9d�FSPD_OVR��a<pC�`�R�COIR�W��N���VF�1l�V�@OV�ESFjP`c�F3f�!�CH8Kh��"LCH2rFuRECOV�T���@�W"pM�P�e�@RO�8�Q�@_h0a0 9@���VER�p���OFS��CN@��WD�Q�d�Q�Q��U�P�TR,� �#@E_�FDOVMB_CiMb�	pB�@BLs"�B+rs!�$V�	���ȩ ucbG,w?XAM�=SpZ mu�b�_M�CpE�ހOӹ`T$C�A�@ހDhR�pHcBK��6�qIO8�q�upсPPA�z���y��u�upҹbDVC_DB��C��1 ��D��b�![�1c��s[�3c��`ă�U��@��QUK�@O�CAB �@7��� �c� fx
��OzpUX�6SUB'CPUr2�@SQ�� sUt��*#�3#Ut��~�Q$HW_C���D@pH�A.c0�_$UNITuTo�>h�ATTRI-P|���@CYCLycNE�CA��SFLTR_2_FI�4�خ�����1LP�K�0�0_�SCTvF_h�F1_r�����FS��Mrm�CHAQ��<�Lr:�;�RSD�`�҅Qؘ3s1p�_TjxPR�O��s0�EM��_�`iST)�:! �)�C!��DI���4R�AILACQ��MFz@LO�P��T7t�`� ���!���sPRE�%S�10�C7���=	�cFUNC�R�"RIN� s�2�Ġ:�f/�RAK�� �ppc�p�tc�WAR�3F�pBL|y���A��������DAsPd�θ����LD���P���do1m��!��TI�"��xac0$��RIYA���AF�P�Aä`GŶ[S�ʓ�MOIs�vDF_���Jc��C@LMOsF�A��HRDY�ORG��H]�v2�ְ>��MULSE��-ST�L!��J�ZJ�R�g	kFAN_AL�MLV,��WRN�HARD`в����� ��n�2$SHADOW`�0��A�MU_�`�6AU� R�.�F�TO_SBR 9��յ@��h�9�B���_MPINFa0~�x�������p��`|A�  d�m$!�$�� xB|bA}@�� �2S�EG� �C�P%�AR�@���U201躰?UwAXE�GROB�F�W��fQ_t�SSY�rP_�hP��S��WR�I��8�*!G�ST�R�E��gP�PEj�HK@A�oҽ B���a���!�P�pOTOr��K@�`ARYn3`+�䡘�UA�AFIHP~�C$LINK���~1K�/!_��at@��!r�XYZ:�:}�5��OFF�`J�)r�f�/�B�@/�����a��3���FI@����:1�R�T/��D_J�AIB�RW�e�0���S�TB!��2YC��.VDU�b?�.��TUR�XÒ�9��X���pAFL�0 g`ǃ2� ����8��R�a 1�K@K�@M�4?�9����"��cORQ���Ai���3H� EP�0���!�`-S�ATrOVE|�2M��1�Ӗ�� ��IГO��j� �E4��H��1}�@ �d��1�}�%�Ә%��AER�Am�	B��E��1@�]$A!c0��[���7�ձ҆ձAX�cIBձ��Q� L�%���)���)���* ���*�P�*���*� �*�*1H��&���)\0 �)\0�)\0�)\0�)\0 9\09\0/9\0?9\1�P9DEBU@�$�;�Gӯ� A�bn�AB�է�q�Qv[@Ġ�r
 Bl�7!CEb�OG�OG ��OG��OG�QOG��OG �OGM�^ G����LAB��A<�I�GGRO��A@��pB_��D&���S�����F,QB(U��4VAND� ��R$��w�U!��qW �q��v�XƱ�X̴�v�NT'�� �
�ERVE�P��� $��g�Axa!�PPO�b��p%��Q��S_MRA�� �d ԰T�`xdEcRREsC�TY.����I�pV��#2aTOQ�$�Lc�$���Ee�T�C� �� px ,P�d��_�V1^2�!�d���d2B�k2�f�QW�� �@@�Q�s$W���fke5V����$����w��"jeOCƱ���  kCOU�NT�� �QHE�LL_CFG��� 5 B_B�AScRSR A)B��#�i�Sj���cp1�U%bq2�z3��z4�z5�z6�z7r�z8�wVqROO����pݐu�NL��dAqB�S͠dpACK,FINpT�4��e�8��.��_PUՓC��OU�SP��guܡ�Dr�v��чTPFWD_KAR7ac aRE�T��PG�ܱ��QUEm���}���A�c�I�/CCss�ڣp?�v�at�SEMR�`	�b���<�.PTY%�3SO�!DDI1���p�Cс�'u�_TM�PN"�NRQb�s�Eߐ� C$KEYSWITCHڣ��D�ڄ{HE��BEAT����E5�LE6b�����U��F����SI�D_O_HOME�OO�7REF]PR��"(����2�CԐO��`�qaO�P3@�&�IO�CM_�YA�SDsH�K�� Dp�o�R'ESUbςM����<ooFORCs�ʳ� ibDsOM6� �� @
D=Â�U���P4�1֦�4�3�֦4�
@qNPXw_ASKr� 0qp�ADD{�Z�$S{IZa$VA2P\�u��TIP��
۠A���``_��H���]�S�C�C2`�y�FRIF��pS0��˩�i�NFe�
��dp�� xx SI�ObTE�P�SG%LѱTY� &���x�C��ҰSTMT�2�P!���BW}Ӵ�SHOWř��S�V����� �	aA00vTT�ߠ\�@�\��\���\�5Z�U6Z�7Z�8Z�9Z�AZ�W�\�ʠ\��A]ƀ��\���_�O0�f�1�s�1��1��1��1���1��1��1��1���1��1��1�1�1�G���f����� �ɉ��ؚ�Q �ش�� T����2��2��2��2�2�2�V��f�3s�3��3��3���3��3��3��3���3��3��3��3��3�3�4��4�f�4s�4��4��4���4��4��4��4���4��4��4��4��4�4�5��5�f�5s�5��5��5���5��5��5��5���5��5��5��5��5�5�6��6�f�6s�6��6��6���6��6��6��6���6��6��6��6��6�6�7��7�f�7s�7��7��7���7��7��7��7���7��7��7�7��7�7�@qV�P��UPDJ�� ��`� {r�aYSL}OKr� � #� i�f����S �4�R@U5;���pRz@8F�!ID_Le��h5HIc:I���PLcE_b��4�$	�v�&SA�b� h`~�0E_BLCK����2���8D_CPU �9$��9�c3�?�4�"�P]�R �|`
�PWp�q FAL�A��S�aKC\AUDRUN�ErAJDrAUD����E�AJD�AUD �T�BC�CJ���X -$�ALEN`��D��@?�RA���R� W$PI��F1�A�42WMp]��C4��.�ID� jQ&\GTOR�@>[D�a<0S��LACEB�0Rp�@c0R6`_MA	�pMV�U]W�QTCV�\�Q]WTn��Z�U�ZС KT�a�U]S�aJA�
t$Mdg�J��D�LU)9a]U�A2A�<���`RaKS"PJKefV�K�wa�wa3icJ�0�d{cJJ�cJJ�cAAL{c�`�c�`ʫf4�e5�B�QN1��\�`�[�P.TL'P_���>�}@p�@Is�{ `�0GROUN0��g�B��NFLI�Ca�=pREQUI;RE
�EBUJ��AfY��P2�X��@]vx�A�G�� \m�/APPRipCT��P�
��EN�xCLO��yS_M����y�LU
�AL�� �7�MC�R�P�B�_MG���CF��0$��␉P%�BRK#�N�OLS�%�2�Rc�_CLI%�i�S��Jr�e�P�diP�ciP�ciP�ciP�ciP6��߱���8B�s�u��# fr�B�A ��A�PATH
�#���#��H�N�xp�`CN�CAt�i��r�IN�BUC-P1y�-C�PUM��YPl���l1E�@���@���`~o�PAYLOAa��J2L� R_ANx��LG@��ߙ���$�R_F2LSHR��%�LO�x�)����7���ACRL_@�v�i�r�ה�BHA0ζR$H$���FL�EX�s�AJ�E� :�O�F]Pȧ�ߤ�O�A]P�O�O\F1ߡ-�A�_)_;_M___q_q�E{_�_�_�_ �_�_�_�_oH�e�g $cedU�w�,o>oPoޡWjT��F�Xl�bce ����ne��zo�o�o �`�e�e�e�e�o�o�o�y���!t� �� -?Q��� A�TZ�eq`ELȰ �*�lxJS��spJ�EP�CTRr�U�T�Nv�F(�]wHAN/D_VB���M0n�� $��F2$�X�sb�<2SWq���v�� $$M��R>���O������厂�Ao0ܐ�n1D$��A.�10@�AN�AA]�/�/��0@�DN��D]�P=�G]@��S�TB���O���N`�DYt@�p$��7��}� �ߡ�:�ޗeg�����d�P������Å̅�Յޅ�T_���� �ത����q��ASYMM���fpM��`h�:�m�_SHrw���{��� ������џ�Jꜛ�������g�_VI����s	 V_UCNI/�$?�'�Jfe 6"d6":�:$Q�G$k& Z�`m���|����%��I����{큕pHH@f�rݙ��!EN��
�DI]���O48�� !s� O�>�I!A��Q�819@�3�F3�08�@;A�1� �� ��ME��Г�a2�"�1T� PT@q��8��1pt�p���8�1�9T�q� $DUMMY}1G�$PS_X��RF�  8��66!ALA#pYP���2��3$GLB_T ��5E�01�@��Y�'1� X�p]w�SuT��spSBRM��M21_VbT$_SV_ER�OWpL_CwCCL3@_BAɰ�O;2� GL  EW�$q� 4+p�1$Y�Z�W�C[`$�B��Ab0����AU�E�� ��N�@v0Ew$GIi�}$�A� �@�C�@$q� qL+p�Fr}$Fr^WNEAR��N_�yFLY��TANC_�ν�JOG?��� ��\0$JOIN�T�!q��EMSET$q�  �I3Tʱ���SM�U��$q��n��MOU��?�spLOCK_FO9����0BGLV\�G�L�XTEST_X9M�p�QEMP�P���b1B�P$US~1�@� 2�sp�C@a��b���P@a�aAC�EpSa` $KA�R�M3TPDRqA�@~duQVEC𠬏fyPIU@a�EaH=E�PTOOL!��c�V �RE�`IS3���d6ÁU�ACH�PS���aO[��3�4�2�PSI�r � @$RAIL__BOXE�!spoROBOd?�aA?HOWWAR��0q<�0�aROLM�2Vu ���dgr��p�T�a���_�DOU�R� H R^cI2���P$PIPfN ���br�ag�@a�p�C���OH0 � D�pGLOBA�6��P����3@�r8�S;YS�ADR7�� �0TCH�� � ,��EN�"1A
�Q_�Dp����R���PVWVAd1� � �`�B5P�REV_RTq�$EDIT��VSHWR��KFԀ��
�A�Ds0
���HEAD�� �����KE�A�0CPwSPD�JMP_��L 5��R��#4��e�I`S7�C�}�NE�`8�s�TISCK!�+M5���F�HNAA� @p�pc���$�_GP���v&@STYj��aL�O3A������� t 
��Gv�%�$���D=K@S�!$,!� x1E50F9P��SQUx`�<B�TERC�0��w�TS��� �&A�W@�ר���x��aT�O�0�3c�IZD�AE=�1PROC�2Ѣ�1�pPU#!�_DYOQRo�XS�PK 6�AXI �zsEaUR�ɳ8�7p��.����_�`@�ETA�P��R����F�
�t�R���l ����ꔵ�榹� ����� ���0�ڵR� ڵb�ڵr��͟��@*��
��s��C)��k}����SSC�@ � h�@D1S��a�0SP20�AT`��⡠�o�~�2ADDRES�c=B��SHIF��7`�_2CH7�*�I�:@X��TXSCR�EE����T�INA�CPk��Dp��B��C@� TU� z@Ţ8�yAV@���7�8��Լ�RRO; fP`7����W5rPUE$4G� �� Y��0S�A�8�RSM���UN�EXk� 6"�� S_ �CB�%2�E�`�%B��C�R�� 1�t�UE{��,2�B��ѠGMT~ L�!��f@O�V�$$C�LA<� �������0������VI�RTU� ����AB�S����1 ��� < ��;�M�_�q� �������������� %7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?^;���AXL�������+�  �p4IN�y?�1o4��_EXEr�8�0�6_UP���1#���LARM�"�OVoP��2l4L�M_P���d^?BOTO fOxO�J0O�O�O�O�O�M, 
6�_j6�NGTOL  �#�	 A   �L_^[�PPLICf��?��0�P�Handl�ingTool ��U 
V8.1�0P/11  ~S-C�(
ya�SW�R^pԄ�Q
F0�Q�U����^p
1232��TOh��X��Z��`��7DC�1�P\�SNone�  EL@T�FRA_ 4��YWbl�PpQ��TI�V�5�S�3�cUTEO�� A�4�9P1�GAPON��n���`OUPL�p1I� �`&tg9�`UB� 1K) ��0x0|0|�����s�1�s����� ��Uvt�H_ur�zHTTHKY���cu� ���#�}�G�Y�k� ��������ŏ׏��� ��y�C�U�g����� ������ӟ���	�� u�?�Q�c��������� ��ϯ����q�;� M�_�}���������˿ ݿ���m�7�I�[� y�ϑϣϵ������� ���i�3�E�W�u�{� �ߟ߱���������� e�/�A�S�q�w��� ����������a�+� =�O�m�s��������� ������]'9K io������ ��Y#5Gek��|BuTO6P�o�cDO_CLEAN�o|@t#NM  ;[_Q/c/u/�/�/4�_DSPDRYRL/?uHI�`/-@@/ ??+?=?O?a?s?�?��?�?�?�?�?<xMA�XrP����g�1X���Q�b�Q�bPLU�GG�`��c�ePRUC� B- �+�/��?WBO\B�/@tSEGF�`K�O�G�A-/ ?/__+_=_O_�O�ALAP�/�N�s�_�_ �_�_�_�_o!o3oEo�Woio{o�cTOTA�LFHI�cUSENU�@�k ��o��BpRG_STRI�NG 1�k
��M�`S}j�
q_ITEM1v  n}m6HZ l~������ �� �2�D�V�h�z����I/O S�IGNALu�Tryout M�odeuInp�̀Simulat{edqOutތOVERR� � = 100rIn cycl҅�qProg A�bor�qȄS�tatuss	H�eartbeat�wMH Fauyl\�e�Alero� ��������ß՟���8��/� �{ �(2���������ȯ گ����"�4�F�X��j�|�������ĿF�WOR�@{��p�ֿ$� 6�H�Z�l�~ϐϢϴ� ��������� �2�D�8V�h�z�PO{P� ��ˉ���������� �/�A�S�e�w��� �������������DEV��D��1�k� }��������������� 1CUgy�����PALT \����"4F Xj|����� ��//0/B/T/�GRI@{�! f/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?z/�`R\�0A �/
OXOjO|O�O�O�O �O�O�O�O__0_B_�T_f_x_�_�_OPREG��PHO�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
.�@���$ARG_���D ?	�����q� � 	$��	+[�x]�w����y�vpSBN_CON?FIG �{ց�Ղ�qCII_SAVE  ����q�rvpTCEL�LSETUP ��z%  OME�_IO����%M�OV_H9�L�R�R�EP3L��pvUTOoBACK$��}�FRA:\��[ ���V�'�`:��W� {� �� �x �]>�P�}�t��������������� )�;��UΟg�y����� ����L����	��-� ?�Q�ܯu��������� ϿZ����)�;�M�_�>A��dωϛϭ�p�����ϲ�INI� ��T�u��MESSAG����p>�ODE_D>���͆9�OF�H߶�PA�US��!��{ ((O�r�߲ۜ� ����������*�,� >�t�b������{�~��TSK  ��x��Ϲ�UPDT?���d5�U�XSCRDCFG 1�v_������|��������� �����e�0BT fx����������rs��G�ROUN)�i�UU�P_NAf��{	���R_ED�1�
L�� 
 �%�-BCKEDTA-Cz���[��P�����Z�r��xW��r/  ��_%A2h/y�F/�/<"��t %�/�/C/U/�/y/a#34?�/�?�/�.]?�? ?!?�?E?a#4 Op? MO�?�.)O�O�?�?�OOa#5�O<O_`O�.��O`_�O�OO_�Oa#6 �__�_,_�.�_,os_�_o�_a#7do�_�o �_�.�o�o?oQo�ouoBa#80�}h�-�Y��Aa#9�lI�4��-%���`����a!CRg/ �o�&��m�Z������I�׏U�NO_D�ELasGE_U�NUSE_qLA�L_OUT ���>#tWD_AB�OR��T�IT_R_RTN׀l��NONS���.�1�CE_RIA�_I)�5�y�FFF���.���_PARAMGPw 1�����?
��.��Cp�  O��Q��Q���Q��Q��Q��Q���Q��Q��Q��Q���Q��Q��  D���I�p����y�����둴� D���Ѱ��"Ѱ*j��1Ѱ9��@�.�?�y�HE��ON�FIG#���G_P_RI 1���� �$��S�e�wωϛϭ�ܿ���CHK��1�5� ,5��� %�7�I�[�m�ߑߣ� �����������!�3�E���OF��찫t�CO_MORGR/P 2֬ h����� 	 �������������̣������q?����p�`�R:Kh�:��Pa�������a�A-��������.
��
��r�@����.��`MCPDB�c����9)c?pmidbgN��� �:��s�t����p�����U�^ �^ ����-���t��0�v����ᐋEgf�����f�/��</� mc:,/T/�kDEF �"(�)@ cebuf.tx��/�
\a/}�_MC��u ԰ d�%�#����-���!5Cz�  BH�B����B�H'B�`�C�B�r�-CZ���D�36C�G�C���D@OC��kD�w�Z=�E��E�O�E��\E�d�E��	F��	?�����%4����<	j���4~j������̓�Ax���C\,Q�DDi�D@Z>�N@ DE�D� � F�E��oF`/R�> ��JBEL@Gb��FO�\G�L��:��  >�33 �����;  n��;�5Y�E��; �Aa�=L��<#׽2i�E�O/��"RSMOFST� .���)T1���DE �� e��
�Aj�;��B��O�O�.TESTRy"._v�R��g��_%6C4�@����� A�A62��;0B�l�;0C(@@c���j�:d�
�QI_����]�QT��FPROG %,�8��o�UT_IܑZ@�䖏��dKEY_TOBL  6��
A�� 	�
�� !�"#$%&'()�*+,-./01�23456789�:;<=>?@A�BCy GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~���������������������������������������������������������������������������q���͓���������������������������������耇�����������������������z`L|��kp�z`ݐ�STA"��T_AU�T��Oe��V>�INDT_ENB+�b��ROQI�;�T2���t�a�n���XCˣ �2�j��8
S�ONY XC-5�6�_	B�u��@�����  ( �А��HR5!0
���+�7=�O�Aff[��o��ß �����՟�0�� T�f�A�����w���үp�����f,TRL|`gLET��� w��T_SCREEN� ,�kc�sc��U��MME�NU 1u <*�o������ �Sǿ�&����\� 3�Eϒ�i�{ϡ��ϱ� �������F��/�U� ��e�w��ߛ߭����� ��	�B��+�x�O�a� �����������,� ��b�9�K�q����� ������������% ^5G�k}�� ����H1 ~Ug����� ��2/	//A/z/Q/�c/�/�)k�_MAN�UALÏF�DBC�Oe�RIG4�5�DBNUMLIM���:�d�UY`DBP�XWORK 1 fk�_[?m??�?�?��]DBTB_)� !�_�Q�PK4�!__AWAY�#:�/GCP �R=|P�6�_AL0-��2�"Y�6��P�(_DBGW 1"ZY�I�,��K?�O�SrO�O�8_M�d�I)PL@+`�COoNTIM3���T���F?I
�eTCM?OTNEND�oSD�RECORD 1�(fk ��O�SG�O�Qm_�[B�_ �_�_�_xX�_o_4o �_Xojo|oo)o�o!o �oEo�o0�oT �ox�o����A �e��>�P�b�t� ������+����� ���:���E�͏���� ����'�ܟK�՟o�$� 6�H�Z�ɟ~�i�w�����@eserved� for Tool �����m�"����X��@mmy $�0E0u� #33 Y������ƿ��������@	! TP K�ey2 (ABOR�@$�6�HϷ�l�ۿ�e��� Pq�5u�9 گ����X���ώ��C��At Rele/ase)q�8u�E��|ߎ����JTOLEoRENC DB�IB�@L��� CSS�_DEVICE �1)�9   �6��)�;�M�_�q�������C��LS 1*����������!�3�E�W�����PA�RAM +`I�i����_CFG �,`Ki�dM�C:\��L%04�d.CSVh�� cd��i�A��CH z� �Oi�Q����'�2�!~l@0��JPѦ�RC_�OUT -�;�m@k���SGN �.�5?R��\��16-MAR-�22 15:01���?1� 4�4:4�5��� Tn�u�-)i�*�o���Im��P��uG�=��VERSION �
V3.1.j��� EFLOGIC� 1/�; 	��(@0����PROG_ENB!O\FR�ULS�G �6=�_ACC6(A��.C�7#WRSTJN�@�&?R�#DEMO,(A0E{!INI� 0�:�5?1� v&OPT_S�L ?	�&�"
 	R575i�V� 74�)6�(7�')5j�2182�$��6?��$TO  ��-@�?�V� DE�Xd'd?U�3PA�TH A�
A�\�?�?O�KIAG_GRP 25���� �	 E�  F,D FAD�`QC��@IC@��nOLkA��ЗO�N�CeECl^O�CkI$C���C� B�m��If362 �67890123�45�B�'  ��cPA���A��=qA�A��33A�z�A���A��RA�A�P���HJPj!@\@p	 ,GQ��A��������B4L��D�(j!
�R�P�{A�P�P؜P�P��G�Aď\A�?�A�Q�*?_@Q_cT�*�б)�^�PUϸP�P� P��P���P��A�ffA�P#P�_�_�_��_o�X_�PZ@`U��PO�
AJPD�P>$P8P2@`,��lWoio{o�o�]`�W�A[�PV�PPP�K
=AE�A}?P8��A2�P+�
�o�o�o��X��`�$PLpx�PqPj$Pc P\�Q�ATPL�� bt����TC@R��Q3a�aKq�p^M=�{G�z�>8Q솅�^M8��b��7��Ŭ��^M@ʏ\Nʆ�p�օE@[P�Ah	 �C@<�C��<�t�=��P=�hs=��{�P^M;��
.��<#8�[ �?�+ƨC�  <w(�U� 4Ƃw���r����~�
��@
"?fE6���8� �����9�k��0�ʟ�@�f�H�����~�?TCzᾦ;�ʥ^M�{��G�^NcQ�����^Nx��7��C��O�
�@�CkJ=C7��Ck�^M������|����`K
�׿%�ED  E�� ��7D+�	�C��O|7�j!8�?6�������9b�zV��6в�eWZ��2���b�����DkC��蚖��#Ϡ���Ϣ{�����I ACT_CONFI���6������eg� ASTBF/_TTSd'
)B��C#��U���MAqU^ /��MSW���7��_P��OCVI�EWi�8��	 �������*�<� N�I��~������ ��g���� �2�D�V� ��z������������� u�
.@Rd�� ������q *<N`r� �����/&/`8/J/\/n/��RC��	9�5v�!
/|.�/�/��/�/�/#??G?[�S�BL_FAULT� :�*��a1GPGMSK�7t7�0T"A� ;ٵ���MC: �C�O�:|#P��OO1OCOUO gOyO�O�O�O�O�O�O��O	__-_L� �<���1RECP�?�:
�3�_���?�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�oI_���UMP_OPT�IONK�m>qTR��L�q9;uPME|J�.Y_TEM��È�3BK�r�p��ytUNI���MՏq��YN_BR�K <��y8EMGDI_STA�u؂��q�uNC�s1=�� ��o'��|,d�_m��������Ǐ ُ����!�3�E�W� i�{�������ß՟|+ ������[�&�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ���2�  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� �������*�<�N� `�r��������� ����&�8�J�\�n� ���������������� "4FXj|� ������ 0BTfx���� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?��?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_�?f_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<r_ `r������ ���&�8�J�\�n� ��������ȏڏ��� �"�XF�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү���,��,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�z��� ����������
��.� @�R�d�v��������� ������*<N `r������ �&8J\n �������� /"/4/F/X/j/|/� �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObO�/�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6olOFolo~o �o�o�o�o�o�o�o  2DVhz�� �����
��Ro @�R�d�v��������� Џ����*�<�N� `�r���������̟ޟ ��8�&�8�J�\�n� ��������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ���� 0�B�T�f�xϊϜϮ� ����������,�>� P�b�t߆ߘߪ߼�� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv����� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?� �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_x?f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�oL_&L^ p�������  ��$�6�H�Z�l�~� ������Ə؏���2  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶�������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x����� ����������,�>� P�b�t����������� ����(:L^ p�������  $6HZl~ �������/  /2/D/V/�f/�/�/ �/�/�/�/�/
??.? @?R?d?v?�?�?�?�?��?�?�?I�$EN�ETMODE 1�>r%�     4@�4@<E7OIH@RR�OR_PROG %#J%�LH�OLF�dETABLE  #K|/�O�O�OJ�RRSEV_NU�M 2B  ��-A)PdA_AU�TO_ENB  qPE+CaD_NO>Q� ?#KEA(R�  *��P��P��P��P4P+�P�_�_�_ZTHIS%SLA+@�S[_ALM 1@.#K �LD�\�@+�_;oMo_oqo�o�o�__R`P  �#KQFB�j@TC�P_VER !�#J!�O�o$EXTLOG_REQ�Vs�QY,sSIZ5�'tSTKRyoU��)rTOL  �LADz�R�A 't_BWD�`�pHVܻqDw_DI�q Ar%STDDLAKB�vSTEP��@>�pOP_DOtbA�FDR_GRP s1B#INQd 	�o�r�F@c��[���w��#/�[�7u���� ������c���ɍc�C�?�B��NB�!�Bz�A�O��B�N΍B����Bl��BM���Af��A�YA|��΍ɏ?��*�c�N���r����� � A�8A���>�����D@
? J6��֑Β�v�b��ׄ�EݐF,D :�D��`E���)�D � E�� b�D+�m�C�(�C��=N��B�ƈ��΍o@UUU��UU���ۯ&�8��� E��@���΍OHc�GP)�K�ƽ6�Jk�΍?x�R��:G:�z��9{����΍�����t<����nLA��������KFEAT?URE Cr%�p�JAHan�dlingToo�l � svde�Englis�h Dictio�nary��
!� 4D St��ard�  f�fs��AA Vi�s� Masteyr��� R597��nalog I/�O(�  90 H�S�gle Shi{ft(�R6417��uto Soft�ware Upd�ate  4 R�R��matic �Backupe�4�9���groun�d EditI� � oadiC_amera[�F_��4�t��nrRndsIm���duc���omm@�cali�b UI�� ER�m�Con��@�on�itor��ct\�j3�tr�Rel�iabt���PCV�LData �Acqu=�:���.�svk�iagn�os��X���cfl�xk�ocument;�eweE���'��Ok�ual Ch�eck Safe�ty%� g H5���hanced �Us��Fr���P�C��xt. DI�O 5�fi�� dwef.��end��ErrD�L�����D���s-����rV���� �p��41m�F�CTN Menur��v`���H55���FTP InF�f�acv�  J�J�G��pB�k E�xc��g�� Pa�r�T��Prox�y Sv��  j�616�igh-wSpe��Ski� 6.fd㰎��mmunic��ocns������urm��F�_� R67�\���connec�t 2��04��Iwncr��str��z�FCB��KAR�EL Cmd. ML��ua��J�Uc��Run-Ti��E;nv#�"
c�P�el +��s��S�/W��  ��License��Ӳփ�$�Book�(SyE�m)��!� toMACoROs,��/O3�,{��IF��H����
 81 ��Me�chStop��t�:�z� T "j�M�i�w� ����Mi�x��X����orc�h��odu�wit�ch(���o:҉�.� d -��Owptm� R7*�ܙ��fil��Pi�ck�X�g� O�AD�ulti-�T������v
E�PCM fuYnT�z�90#ow��RegiE��  td���PH�t F*� D/�[Y�Num� Sel6  r�y��y�� Adj�u����k�w� � pr�tatuR*�NDI��ٵ��r��RDM Ro�bot�scov9e�*�Rem4 ��n� ,���	#Se�rvo� ��?S�NPX b��(�r�t �w�Libr���pbo��w��9 E{   m� W �o��tm�ssag� Pv��!z�[s? in VC&,�Ħ��` ���(TmP�"/I�� )��� MILIB=f�xtp� P Firm��)�d���n�'Acc����e�71�TX��L��� eln <I0� ���e\mc�1r�quu�imula|C��� te.f�1�u� Pa���Ma���T��^Ѡ&��e�v.�Ѧ�USB �poo @�iP�a�� ��,@nexOcept��# n�� �\@�����n0�VC!�r���:hk�1<�j4<�{+�4�<�SP CSUI��к��IXC�&r�o�Hx�� 
�Web Pl����97��QC!�N l21R���ԩ�D��3%F�� i�gXGrid~!play o��gX� ��L� �iR^nIVMRe  e�� -2000iB�/165��rAs�cii���1�� �5 (K�UUpl����35�s!��!t� rc��Cyc8t���]ori��5%7FRL��amY*�HMI Dev��c (Y!����PC���-@o #asswo�&�2
49\��64?MB DRA�!	�l2�bFRO�kY�7�;rc�visD���95c���ell[�L�7H54�sh*q�	"�0C|c�^�2@Eub��p�6JDEutyt��s��VIct�� .���� ��sp� 2��aV�B b�y 
 ��	 B"X�q� it2���T1�>�K%.10�OL��`SupB�Rc��OPT ��njN�S �bS�B�cro���c	#{%�T mj�p��='�a�pues�t*�SS�`e�t�ex{� ���$Li3mipYb�Sp����1��0P���gJ�n�Virt��	#����Mdpn�8��h{51>CVIS� �IRpvC�JDIR�CALv>D�+�I�C:;0x ��p�hicD�hо�Ab�ui�l�� F��!PMM�p�� �!flowh1f.�sk�OSFILE� Ar" u�co �gtp��BMON���IX c�җ!m� T�N@PTTB:z��i��R805� ��J����
��⊔�j�^�m����"P�ALT:�`clu�d���AIW�- �Wait/Y�ean�� tk��TP�b�DOES NOT RESTO ��60Lin��mar9k��useJ�z ���c�  Sync�hr@�z���DSU�PPR��PRG _IN AR�A ���Ag��OVC_V�ALUE�OBL�EM ��V��TM.i�TMW��G����ab�A MOTI�ON�STRUC�T l��BRA�KE ABNOR�Mx� ��g�$F�MS_GRV0ISMATCH=uu�Z��MAST HANG UP 37m��MULTI WI�N/LOCB���S�ERVO��AG �GAR*�
�GRI�D DETECT BUA���!0������TRANSLA~Y�OF UTX�|�F DB/s��DO PULSE�@ENCCAME�RAǁ�c�`RE�MARK FORh�� w�L�0\h����EXPANDED POS>����%'����SCRE�El�AY CRU�SH �P!�OTN560����fԡ��ND�SYRUN�NI��Ɛ�US}R��F TOLp��NCE ��vK�F�SE��Ŧ ���S�-144 A��AcRT��
p�FA_�� CPMO-07-3�wAUIs�0��'mpl����ڢ�Cpsᇡ�����R>��sydem�ַ���A��snosv!.�����޷�i����gA S���HQ��aV_cmC�-PH�qT��!  ORs�PA&;6�`�P�R��[qdp�(CQo��Y�P,�" �1 �ҷ��G���ҷ�g�R556�ִ���i�c��e�|��G��t�g��2�G���aHP �spotplug�N�Sp��O�-in�b�SPPG ��0~�r�(SC�P`��qLC���J�\sw'���  ��� t���^� ���trsvy\���1.pc
�\��  fx_�2�����%3��B	4!.:�B��5��D��&6�#�C7�	���B	8���Btn�
�0���=�F�n��s�N�Nomi�p P�osi�Q���NN�549~�Ї��`(B�ѝ���TX�P5
n��os\n�mtp "NMTX" #1�П]�et6�OMP�.����-fxu{ifN�-fle��b�FXUFd�Ё�*"('�6	"$  �f "*!�sq&_ �еo$�	 ,]��t#w��rl�o(u�f.vr.��'�
@in�cusA.��3&#2+1��"�� M?U4K?]?�?�?�?�? �?�?�?�?�?O#OPO GOYO�O}O�O�O�O�O �O�O�O__L_C_U_ �_y_�_�_�_�_�_�_ �_ooHo?oQo~ouo �o�o�o�o�o�o�o D;Mzq����t���� ��	�   7j$���v|��r�q��j847\wti�v��/���a��/�q���weW ��=����47,r76�8R�asyArm�&�fun?�f�C�R� S01h���:��(X�t E�����X'�~�\popupct�#Ã,���aN�M�-She{lld�R533R���J� (Mu��-�[���;'���vrdbc2
5C�%� ��enio.fC�E�nH�ced I/�Od��3���J�6�v�ŗp��ܷ���re�pa��c���?�ac_cuairR�AP�GAirS�6;�0�kz� (\�p���O���S�ca
���4�O�� �2�!S�� 2 �Guc�����49 GR63z����(��P���@��g�aΠcib�#A�oSEL��^�/���!C�`�n>,aflowL�3�� AF-AS-F�MS�mmP�AFSM�x�2~勁����(غ����S�˴��afgl
2��G�@�!��̴ۢF�̳2V�F�e�AFް���@�������᳣�O/�e�2ȡ̱��d�:̱2L�AF2�Ͻ�2�����l��RӋ 1B�sŚ���x���!Aw����G�_�ɶ3��qA�!㹽�AS �� ~�5������`#����v�LO��.����˱�ݻ��C�clr�pthR�ic �Cl[���thϜ7+78��7��gv�ȀBas��@�����  �ᛲ��>�S��㒐���tpe=���s�sub������n��=�� /�w�set�����"��q��w�q�Of�f-line S>vulari6�>��85>���[�85 �( ��tya���s�iad\tp� "SIAD�/�����,k�plu�g��Dispen�se P� j�=�S�PLG. 9s�(���g-i��� ����ea�\sld�spi�"�U8���0�� L% Trk F��̀<��>���p�%���For���tq���(�]tcyc "T�����k�tgtp�/��!�l�la��-#ptkmisc5#�" !����w� ~���osable EOAT<�_�G���@��(@��
� ��3Q!�b��"���%1��Fo�u��os1�)t�4�7
���47 (U4��on�)0�_� K1�2+3��7��a�J5��r70��erv�o Tip Dr3es�08>��"�0ȁH7�r7��~A\turnd @�b���D�'�����M	Hb<+�2	��@_��Lq�32]?C5/�S��Ain`�� ���'ggcht ��VG���r�SGCH J*!J643>�Q��GN CfQ��cT\svsvch���CH/���TglgsouV/�[gnc]���_�P�R�	dV;�s�gdia�Ssb �corey2XDG��P70�P�Q{<�b(�~d7�`O��rc�cin�ib���^btdw�j9�52Ҵut@un�SCS<���R Jp�iH8r({��u`����q�Pat݂ c�w�����ux�h869I�7�wl�

/F,
1�v��3� mtsv? "MTSV�X�j983\R���&P�s�ov��&_p�^��vruk%_c6����� ����pex8_�r�col$Q�����v�v"�r���&�s~xcM.Tool���k��=MTOF�7p84 J571 R814�!7E���(��q���	mtofs�0��ߘ�2�⒑�pt�a��l�leto���k�PT�LC�9����J9�813���H��� T�4�9��`k{;��1�a�\pmk920 "K���S!R����1P�Ȥ<���2¢2�_�ި4���!�ڣ�a
6�1¡4��0�����E�ܣ�q8�4f�4C�c&0�5f�����ݤ��9�7f�7C��ަ�gr@"GRIP�".�쿶��1i "�OPTIC��1ݧp�alf "PAL�F�Q��@�{ĻPS�SUC�F!ަcpt "UNIT�S7mަ{xf�XFER��,ԃ��et��L�U��&ʾŏ��psys�dj��/����mޤopti��Kޥ����7߹�ssu��+�ޤ0cpG!W���er��S�N�t�ߞ�sӸ��d+��[�adpՂzaAd�apt CtrlLF�3q50E�G0���_���l\apIa��.�C����a�1�l"�gui� GU!I��T���c[�c���xogJo^U etra�&��u���86F�� �(���r6��re��3�ETN;���.S�X��5x���j722\cust_wv6�RS�Cv7x�RS�[8��;QU	9�KUwv�102oRwvpa�t-�T�ang�e/;Uh`#C j8�0�WeldCo�ndMo���H�J`K�#7a�Dq (T����iJ\atk3�0e���R�1�{�w�m]MON�_�0\�$�_��$Xg���p��b��"Atx��%stop�/�rù���Zd��y8�N4Cir��ld Pr��XvF�ׁ��K��1��cS7�OF1�1\q�-\?8�a?t_ufrm.� �#ER�7xcArc �Abnr�l \i�tob9  ?H552}�1�21 [prc��2 a�1A�AVM ��20 ~��J614���@TUP mch� "#@545�P�C#B6��VCAM awam�0�CRIMe_@UI�F��#A28 0`v�r_@NRE�b.@R�631�s�0SCH���DOCV �lisi
@DCS�UE�#A045pR51EIOCe \t��0542}�R�A�96 pC
@ES�ET ��c
@J5�K@��#@7K@;b�MASK acr�yv@PRXY c�w1wB7%��0OCO- Pht�B3�s;B�2  Q�B0�p �pa#A@4�;A39��0Fo�@H^SI��LCHK�@59>�@OPLG ��;A�03 ��PHCR� :�PCSP  �GW�R6 ��;A5�4��PDSW@_�f�0MD;P "F�O�@OP;P�PP�RO!ÏB7 mf�ork�B0�UPC�MF	e�@4f50	7�U�@5-hg��!f�RST-f69`c;lmPFRD@�S�RMCN	eH93�0�eSNBA�US�HLB	eSM�`m�exte�B6�fP�VC-g2�`��~QT{CP�UTMIL	fw7895@ups�`wPAC�fPTX	e�TELNrd�R9�Ef8@w1 mpwush#@958Ef�957	eUECK�YuUFR�fVCC�M	eVCOR	�k;.vS@IPLU�@�I ��_f�qXC� kZ�_@VVF ��WEBP lY��aTP��t.�p�R626 T I�npCG�pnF��I=� ��6�P�GS�R3_q95 �718 P�073�8 f��1�@
  À�AC`6�A63� 794�B523n�5R65�1SuaO553 ��A4�@�gC=@1qED064_ tamapF����O�6 sths�._@LIO ��w�^p��5 - He�fPCMSC��ӂP���51@STYLy t�_@TOP ����PR5{@Wave=,�PRSR ��A[801UOL�Ph� v@OPISY0��`&� w.��0L�p}���S��t^pET�S�fun�0SL�MTY0��B9 6�23�A�`E�5FV�RC�0_��NL 9tj�wp001E���2E��3)E��6 j��:@U0'@BDݐ95MEݐ8 a֐��U0�`6������Q5��?@s@S����0F�61�=�3� ��;��@69�U�5`*�faF�_�7� ��݁a�8Y�04B^�9��_�_PT�up"��20w0��6u���c7 ���@��8 �"Z��9u�us�0U�1aw�㢸�{@Ʀ�@Ҧ�33ݧ38`���`�
�@�7 R.$�M��/�K ���9L���40E[�1̀SSe�@]�2��Ea�oANRSل� �334���拰��n�=e��Roboz���net�����ደB�9���!拰j��\srvo���4�@�h��x�����Sr}v��t ROB:P%M'�e�4��5��G��n�r��b*ŋ�ite��ӿ�5�-��̝6��35v��56�4��7@Main>��tatio�����6����������o4�ŋ�S��, '���苰 拰\��\cc~�� "TORC���������L��cr�V�CR�����5>'�xk965���@���N���MО�6��0���;���o_��w5���0ch��y6���Cv.j�k��iw2 ��
��x5�����2.���n���3�V�h�z��5���uSif����c��_�3E@H��,�l�����"T�1���T�2�(�Z�l�4z���?������/�l_i��}3���勰0� |����  �Y2?�jog\dj�ui���og��a�wmfr� f��F� ius�� Eq LibJ��6K�p�S�/3�� (��b,��2�7�_5'�\x���� "MF��(���d5a��n7y57eM�� mK��߽Ҡm���g �����̞Atw1������tw���#���N6 ink��0LR 8.��6��J852���oJ597�98��88�J�!�1^%N6���b�GN ��k\e3tl�@.�CO����O#A` "ALNK8
�>�%rd_�PB8�� �"\wr*1OD=�"lS ��P$d��088����PN wARC��PRM�3���B0��Nŋ��!8x^����1SU P� �$P��Ç�H���0���pм3mpana�/'�ȣ0�1��H57,X��85n���� �ã0K�BH@��<��1�bel������R��<D41��HDY<�dhen��8 <A��D���Cm���EN������D.��Ex�ن!� kemp�ЬD¼3�m:re��2��pEf"sFMImG�A00��37JR���P�!�IGC (�P.�E�%�чߑT� wavs��IGE��>G�migco`'�mn&NA�ц�f�avavtj�VT�Po/lfrm "�S�pGoYmsy�AS�Yqo/lpdhV�P�DH�oYktpdlf7�DL�o/lrf�`CRF�d�y�p8�t3b��s�`.vrb3hy�rLO5ccr� �p�4c�§�Āq������������R��R�Sg�S����.�o���.��Z=fArbt�\�`c.2  ��� _	�b��! Tert=iB
ELS�P�2��Ug��YL (C�ommyle seU�%)��bգ��s��'�ps01 �"PS��.#le?\pscol���ul.т�ry�Pr:� ��vׁ�Q�4syr�sr��-���ic?e Requ��g%N��SRS�2K�9�P�645.�9R S��"|����(����v�b��/�,M�ۂfO� A"��s�O��sr�����aP5A��+�qm���2813�P6�49Z�89�� �A�{��Z�.���g�#st�M�\����p|�
?�M�utl��v�'�&Q�N����q ?spdramj�!�/peed.�pf%�QΊ�NN05���J6A7�2NĻ�� j�(��d RH�-�	D��b "RMTX"���ƏE�  ;�2 "S�0q�pQD���slmt�7oft� mi���SL��H6Q64n�H62F�20��607B��P�38e�2 Hk�e�s�;�m5l�62K�79���795�79��6�09j�1F�1x�4���5��2����H6���843[�2s�8c25j��6�MT+��"���6����f� "����S���\f봆봖�0n��- Positkio�l��esf �봷1N1h�ݻP(,���ti��,봥��ǀņn1Z�PO)Ss� �0� ��h873�r�rive Axes+˳H8��4di��(Dual Dr봑sΕ�Ȅp��C�\�B�j�.�kŔ*�e9x�sj� De)��1�63����AM? Indexjź����&�\ami0:�s� �mi&�8��ca�sC��nt �Angle+�CO�;����봗#COM��Mom����������gou���!� ��
fl���Envi� m���6kŎd�820)����f�l(�2� |�r��ionΓ{�ǅ�K�r772\ic���$	� �x0Z�˱;��2atznȺ����c�TJ�yn�cIns�p��R76�� �#���Xj�GrmSB����T�zb5mK�masyA`�jբ�nc\��MASIr�{���bas��ultiC-A�`�6V��7v!0� +��5k�NN�P F��se��!\��FRLK��v�k��hdzՎF봅"f'rlk��&�m
ŊTir���C��il/�-&e��r7��0Zond ��:����? "ICRZp�%�Qg8�Piabic�.T�IAB0c���0o�e�I�0V�0E �0��1 (�1�4���0濡�0�C�2\5i�0t� IA˱�p���"�@AiciA�C�0b��!�1�1��!ޛ0main�sDP�1n C7`[��0e�DLPV�2�0��:hpV��P M_@��@̘��O]B�ưI:A��Єdp�CD�(O�F"�0N>I�A �B��0_�Fd%4��eo@nn Sta�n�A[�'"� MC�N�>�90�096:�s�5j��0�Q=����H�0���Q�2~Q(R�em^PkAeSdar�dI0��W2�NQ�0\�tprcmuǰC�MU�ku�1�TRP\rc�0�q��jBRSUF�173 �0uipp��[��Ae�J61S �59Q�I�0taV"i Eq[A��Ζ�Rǅd�!ȡjt`�Pcp�����Esr��A�Qvb2� �Q⦷ka�@xa �0#�-���1 �a:���1 awmgenyl�q�0ener���Weld zQib�oX�0AWMG�U7{o _q(G>t�A�`%�b�;�d�60t[A3r�t�1.y�R msh�cq@�3��n sh�e�qqGR��1CMSC�U�A���RhjQ�(���p�0l�0rd$�1F�8 p[a��u\q�sh� PSH���� X  ������0   ;(L r wKq�1K/Fe$�Q7�Ij��w\cl
A "J�����0 H\j�Qcle��"E�S�HeӄuybU��`{A�ybmdprm"�8�zali_varsS�<���iconu���dbg"��0Iz�ց?rgpged"��1l�&��� Ԅm_�0�1�i�Q҃m102<؟�e_no��ȕ�wrspq����wrpirS�[q>��0�gas��Y��1��_�s���wr������fyfӯE�inch30|U���extwd����wrc����'�DՂrdS�Q�D�0!�i�����aN� b�i����0�Ə(��/i��RF�p
q���sa�j�ca��ntKCM'AP ���O D�B��)�T�f�ap"Qj�A�PC��Z���0st�m(PSTM.Q{� ���apcevre*a�o��in
Au7a�*a�is
�rbCI�SD G�QMetae/`�3�0T56���i<�cQ��Q7�ar� >�,KQ�Y��(�\+sl(�gr0S�14�e���q�	B..i�A�����d��/�[a��>�@�1��Q�d+Q�G 
�	(5ф�M�Q�O K�� ��`+�2�`KQ����@�B��Kq��GT��sU��0ӛ0S30le Act�C�8R��Y
AQ�4.��1�㵏�IZ��\J�ds��SU ^�%����{A�#���s~�!j691.f�1�ServoTor�ch9��6Jv�K� 91 (�K�A��.�Qsvt��VR���ARC
�es4 F4���Q4��MU�dq�v�z�vt/���5� +QtFEv� ՛0"S`��0h for �Alumi��98�2�� 82�����w� ��	���d�{���oo�q��l���L�ϊ��\srvt.vK�3e��0`�hP�AS`�� A�༫<
�S016F�8P5��0�*�(!ez�0��hS�ATNQ����h
�"P�QNGС�	��2w�ADW����t��ҋ�8��wenmr�8s�nhanced wMir�bmag �n�bR69�Q90�2+�E.'KQ I>!���I""\mjQr�MSIR�c;� � e$!�.b�06b"%�tmbu�stcpy�Mod^�  TCP��RE ˑX nvkAd�8���!fKCP>� \�$��Pm:1"MBUI 2���i2d0� i�+�%ܛ�p�930�sPR�OFINET��O\J���J93+� �0 (�5��>鋁Y�3~�Ppnio ":����x�1"P�q(@RIO�/ǖ$A��u�3)tGj96Od:��@gT�UHc67J�O��Q�`FSW䑡@���?�K67\fswp�r��W+F�}�A\f_�ach޷	�A;b�er4���96�p_�fwd!6���f_�rea/T[O 'Qn#eu4��_�Rr��sR8��C�Qurn����%Senא� $Ss�w�t�_fswcol�#�n�AQ��A>k�cvvcuj�2��iRCalib �Vz!nc Utl�4�VCUT� ��1�?�b(�a��Vis�Fu�cj���`k�vSccU���c�tpfia�_z��`p6bp�_+�apset�3���c\z_�p{����k��uKA4���c��j�988/�To��o�rs1�!�p.�=8j�? �p ^ol �+!��+��p\gf *��D�sT�c���VMas@��9�;� |�����1� �Posij�����o�rdt���v�
�02\��up޶�����r_dc1$AB�A!s.��I[\N�b jAn�e��b���� ����ۿ]���+�ޘ��� _wQW�� k�_c0y�t{G���F4x�1k�nifi3 �speY��94� a�1�UI n���v��>�k1��`�\frc1o��
�j9��1��Brake chB:�f�`0�{Q�5G5J��(�ck�rp�X���˕51��b��BRCHUCD ����(P����5/�C�����mulaneou�s�=���>55`�l�oH�Siɀ�STD u�LANG ��!�cs��0C�T��?\cscsm���1ﳔsﳠ�=��pCﳡ�N�dss' �ﳣ@c S�F��
�����3�V6	8��F�,��sﳥ�s\��u�ߣ�Ĝ��N�r69����gonost�eo� n�����1�U�i-��9��C�ﳵ��7�!�\�"DVM0V����"r6�Đ��! !��p��9Uԧ� tr�D!Dﳆ�2ﳡ�[�4� 1TcԦ���er�!��|q+�\pc3j��p���Ƴ075.�os.Re���rN� ��g��2c�6��ė��� �����75\pt�TJC6���b�� �����Bg�ė@�I>�S�i>��8�0�J979a�0a8 1���(Iep	i{�UL+�oﳔ#��a��f "NR�U��¡�prst�a2�£��gutl�.��RBT��O7PTN�q0\?�r0?V�@H nr?�r0ovq?l rb?rDPN���!�rrdfi����u����bascic�ߡ�fc� �J��A-�q��H829V �$��9�@������P}h�c "F2��
Ӡ29���j8y3��ce C��tour� UPD	T3�5����3Fo��on����a��Ӵ�Q8�hoff���r� 35�fnV���r��\f�V�����\fcn��rg%H3(��% ��r�A �����6�%�D�E�������g0=��$���$n(��/1!46%u��C/ T0\> ])A��av2tp�0ޖ�0v�0��2v6`�0���0?U8 �0�1Br�0���0�4U0>L�vpofs`1|���1�3y0� mgp�s�0Nv�<un�Q�,x�0�4se�5ҌBT0���b cellf�1��el�0Cp��򠄫1��R�1�f�B��5{19�1ll F�B��0��p�0b�C�Bn^�0fncl��"RA���Z�0^V�Bfnd�ru��AsIND"p�1�>�A�1\fn��t�A^f�0t�B&PTPexjA�?�@�0%QTP�c�1�v�1u�B&Ptqd~_�[ Q�2�V�Gj7��0- V�-500i/�010i 3D�0� [S��15�`ab`��13DE��0N��<9\calc@�_.2�7�0vsfit3@Ep�0�{a���07�u��0`�`Tra�0B$��KJ�a�MJ�`�b �e�1�bE��10Ovz�0j�`\que�1�?�3Arpo��8_�`}8�1epush3�#� ���0}s\�М�1v��/�qkm�1ޕ�\�swa�?�h�qa�inj|wkclb*O��?qvs
AJ\udsblt���e�enn�g�|wig�chk��uv�av�uA�s�� �|��0 � �тv��3��_p`��FA��GA"73�1Gcro����,�v�A#po ��0�8�a��jB��iR�qon OErro9���.m�9FQ�A757�Aж<�1�� (iR�A���R.]kZ�<d\m_herhd�AH4Px���}��\ire:AR���ree���/0H�B@���l��Z�h:Ahd��� ������j���cv�a���`�1S?P APAS�A���SASz�09 �q �CTAMڠQTA�BڡP�AGz�13�Ҷ�Π(�`�Q�����p&u/M��pas\�aama�s+�=��
AF��c��s��bia0�B?����VS����VSIAС��D��q����(�A��vAC�  �6�� ����1  !   뱚�� �Ó0(��8 ��\��}�ұ(H� �>�]ia\ia�`�aШ`���P�g�Qoi�Zĳ|c�������  ����*S�YST�EM�0�A ����$�ˢ�S  ���0���������ATSTKS�IZ����/��0���� ��+�=�O�a�s߅� �ߩ߻��������� '�9�K�]�o���� �����������#�5� G�Y�k�}��������� ������1CU gy������ �	-?Qcu �������*��Ȳ��TART�_T SAG���$D��IGNAL���SARTUP_CNfQ/a/s/�/��/�/�/�/�(J�:2!
�
 �/? ?)?;?M?_?q?�?�?��?�?�:99�$�K��$FEA�T_DEMO _C����1@?   �8M O OMODOVO�OzO�O �O�O�O�O�O_
__ I_@_R__v_�_�_�_ �_�_�_oooEo<o No{oro�o�o�o�o�o �oA8Jw n������� ��=�4�F�s�j�|� ������̏֏���� 9�0�B�o�f�x����� ��ȟҟ�����5�,� >�k�b�t�������į ί����1�(�:�g� ^�p���������ʿ�� � �-�$�6�c�Z�l� �ϐϢϼ��������� )� �2�_�V�hߕߌ� �߸���������%�� .�[�R�d����� ��������!��*�W� N�`������������� ����&SJ\ �������� "OFX�| ������// /K/B/T/�/x/�/�/ �/�/�/�/???G? >?P?}?t?�?�?�?�? �?�?OOOCO:OLO yOpO�O�O�O�O�O�O 	_ __?_6_H_u_l_ ~_�_�_�_�_�_o�_ o;o2oDoqohozo�o �o�o�o�o�o
7 .@mdv��� �����3�*�<� i�`�r�����Ï��̏ �����/�&�8�e�\� n���������ȟ��� ��+�"�4�a�X�j��� ������į����'� �0�]�T�f������� ��������#��,� Y�P�b�|φϳϪϼ� ��������(�U�L� ^�x߂߯ߦ߸����� ����$�Q�H�Z�t� ~����������� � �M�D�V�p�z��� ����������
 I@Rlv��� ���E< Nhr����� �///A/8/J/d/ n/�/�/�/�/�/�/? �/?=?4?F?`?j?�? �?�?�?�?�?O�?O 9O0OBO\OfO�O�O�O �O�O�O�O�O_5_,_ >_X_b_�_�_�_�_�_ �_�_�_o1o(o:oTo ^o�o�o�o�o�o�o�o �o -$6PZ� ~������� )� �2�L�V���z��� ��������%�� .�H�R��v������� ������!��*�D� N�{�r���������� ޯ���&�@�J�w� n����������ڿ� ��"�<�F�s�j�|� �Ϡϲ��������� �8�B�o�f�xߥߜ� �����������4� >�k�b�t������ �������0�:�g� ^�p������������� 	 ,6cZl ������� (2_Vh�� ����/�
/$/ ./[/R/d/�/�/�/�/ �/�/�/�/? ?*?W? N?`?�?�?�?�?�?�? �?�?OO&OSOJO\O �O�O�O�O�O�O�O�O �O_"_O_F_X_�_|_ �_�_�_�_�_�_�_o oKoBoTo�oxo�o�o �o�o�o�o�oG >P}t���� �����C�:�L� y�p����������܏ ���?�6�H�u�l� ~��������؟�� �;�2�D�q�h�z��� ����ݯԯ� �
�7� .�@�m�d�v��������ٿп��   ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� ����������
��.� @�R�d�v����� ��������*�<�N� `�r������������� ��&8J\n �������� "4FXj|� ������// 0/B/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�? �?�?OO(O:OLO^O pO�O�O�O�O�O�O�O  __$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv���� �����*�<�N� `�r���������̏ޏ ����&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ���*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?|?�?��?�?�?�?�?�9  �8�1O(O:O LO^OpO�O�O�O�O�O �O�O __$_6_H_Z_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�o�o�o�o�o
 .@Rdv�� �������*� <�N�`�r��������� ̏ޏ����&�8�J� \�n���������ȟڟ ����"�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�?P�?�?�?A@�8 O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ� ����0�B�T�f�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r�������຿̿޿���$F�EAT_DEMO�IN  Ā�2�����IND�EX'�6���I�LECOMP �D���h��5��^�SETU�P2 Eh�~r��  N ���[�_AP2BCK� 1Fh�  #�)�����%�����k���/����[� ���ߌߵ�D���h� ����3���W�i��� ������R���v�� ���A���e������ *���N��������� =O��s�&� �\��'�K �o��4�� j��#/�0/Y/� }//�/�/B/�/f/�/ ?�/1?�/U?g?�/�? ?�?>?�?�?t?	O�? -O?O�?cO�?�O�O(O �OLO�O�O�O_�O;_ �OH_q_ _�_$_�_�_ Z_�_~_o%o�_Io�_ mooo�o2o�oVo�o��owɫ�P�� 2>��*.VRN�`*Qw�c}���e8pPC���`OFR6:��~�"��{TF�F�X��uC����)�����f*.F;ُ�a	�sǏ����*���STM @J�S�^��pK����`�iPendant Panel����H���p�ϟ���3���GIF=�g�r��S��"�����JPG ���r�ׯ����;��z#JSE�n��`�\���%
JavaS�cript��ůC�S���q�߿�� %�Cascadi�ng Style Sheets���`
ARGNAMOE.DTMϰlu��\a�ρ��Ģ�N�	?PANEL1����%u���%ߜ�����2߀��n�+�=�����3�����߯���V���4"���v�3��E���Y�TPEIN�S.XML��}�:�\�����Cust�om Toolb�ar6��hPAS�SWORD��n�FRS:\y�8� �%Passwo�rd Config���o����9�o ]����"�F� �|�5��k ����T�x //�C/�g/y// �/,/�/P/b/�/�/? �/?Q?�/u??�?�? :?�?^?�?O�?)O�? MO�?�?�OO�O6O�O �OlO_�O%_7_�O[_ �O_�_ _�_D_�_h_ z_o�_3o�_,oio�_ �oo�o�oRo�ovo �oA�oe�o� *�N����� =�O��s������8� ͏\�񏀏��'���K� ڏD������4�ɟ۟ j�����#�5�ğY�� }�����B�ׯf�Я ���1���U�g����� �����P��t�	Ϙ� ��?�οc��\ϙ�(� ��L����ς�ߦ�;� M���q� ߕ�$�6��� Z���~���%��I��� m����2�����h� ���!�����W���{� 
�t���@���d��� ��/��Se����<N���$F�ILE_DGBCK 1F��� ��� �( �)
SUMMARY.DG���MD:!a�� Diag S?ummarybo
�
CONSLOG�W:L��tC�onsole l�og�n	TPA'CCN�@/%(/e/�pTP Acc?ountin/o
�FR6:IPKDMP.ZIP�/
�/�/q� Exception�/��+MMEMCHECCK[/�Pq?��Memory D�atar?ra,]�)]1HADOW�g?L?^?�?�3Sh�adow Cha�nges�?�-��)	FTP��MO�?QO|7�mment TBDzO�r=t)ET?HERNEToO��01�O�OtEth�ernet �figura?udA?DCSVRFnOTO�fO_�1%DP �verify a�ll�_�10"�?UDIFFw_]_o_�o�0%�Xdi�ffo�W01DPCH�GD1�_�_�_�oc o�o�S!�Gi�2ofoxo 8�o4�oGD3�o�o� #�Gv�UPDATES�.�p��FRS�:\��uUp�dates Li�st��PSRB?WLD.CME����Y���PS_ROBOWEL�O mޏ�����8�J� ُn�����!���ȟW� �{���"���F�՟j� |����/�į֯e��� ������T��x�� ����=�ҿa���ϗ� ,ϻ�P�b���Ϫ� 9ϣ���o�ߓ��:� ��^��ςߔ�#߸�G� ����}���6���/� l��ߐ�����U��� y�� ���D���h�z� 	���-���Q������� ��-R��v� �;�_��* �N�G��7 ��m/�&/8/� \/��/�/!/�/E/�/ i/�/?�/4?�/E?j? �/�??�?�?S?�?w? OO�?BO�?fO�?_O �O+O�OOO�O�O�O_ �O>_P_�Ot__�_�_�  �$FILE�_�PR�����P�����XMDONLY� 1F�U�P 
 �;_o__6o�_ Colo5_�oo�o�oUo �oyo �oD�oh z	�-�Q�� ���@�R��v�� ����;�Џ_����� *���N�ݏ[������ 7�̟ޟm����&�8� ǟ\�럀���!���E��گi����ZVIS�BCK�X�Q�S*�.VD�a�ϠF�R:\0�ION\�DATA\L���ϠVision� VD file ����տ������/� ��@�e�����ϭϿ� N���r�ߖϨ�=��� a�s�.ߗ�&߻�J��� �߀���9�K���o� �ߓ�"�4���X����� ��#���G���X�}�� ��0�����f���������U�ZMR2_�GRP 1G�[��C4  B�> 	 �Q��� E�� E�@����`
� OHcG�P�K��^�Jk��?� x`� :G:�<�9{��H�A��  dvBH�C���N�B�ƈԜ`�� z  D���>��	o@UUU�UU��`/���#@=�udѽ��H=���=�~�=��yC,���;��.;!�9����:�b:�l?��/ /�/�/��E�  F,D] �!D�`�#�u��-��E�� �!D�+�2C�dR_�CFG H�[T �/O?a?s?��NO �X��
F0�1 �0 ��  �0��PR�M_CHKTYP  �P�> �P�P��P��1OM�0_MsIN�0<���0v�PX�PSSB%3]I�U�P��#O:CCOUO�UTP_DEF_OW�P�:�YpAIRCO�M�0{O�$GENOVRD_DO�6��R�LTHR�6 �d�Ed�D_ENB��O �@RAVCrxJGC� �� [OF_�/j_�x_�_l7�P�QOU{ P��B�8�(�_�_�_�oo  C�f`\�Vo�X�oYm%~oB����b�	�Y\OPSM�TSQY� @ed��$HOSTC%21=R9��G� k M:}k;�8  27.0z�p1t  ek �����z��1��C�U�x|�	�	anonymous|� ����Ώ��7:� ����ik�P��t��� ������������ 9�ӟ��^�p������� ����+�-��a�6� H�Z�l�~�͟����ƿ ؿ��K��2�D�V� hϷ�ɯۯ����#� ��
��.�@ߏ�d�v� �ߚ߬�������� �*�yϋϝϯϱ�{� �Ϻ��������Q�&� 8�J�\�n������߶� ������;�M�_�q�F ����|����� ��0S���� x�����K!3 /Gi/P/b/t/�/ ��/�/�/�/�//S e:?L?^?p?�?�� ��?	?�?=/O$O6O HO�/lO~O�O�O�O�? YO'?�O_ _2_D_�b~qENT 1S�[� P!�O�_�R w_�_�_�_�_�_�_  o�_,ooUozo=o�o ao�o�o�o�o
�o�o @d'�K�o �����*��N� �G���s���k�̏�� ������׏%�J��n� 1���U���y�ڟ������ӟ4���X��QUICC0e�A�S���w�1�������w��2���T�!ROUTERU�1�C����!PCJOG�����!192�.168.0.1�0~�s�CAMPRYT��ѿ!�1���RTn� �2ϓ��YTNAME !~fZ!ROBO����S_CFG 1�RfY ��Auto-st�arted�4FTP�?,��?�OW� �?{ߍߟ߱���hO�� ����@�.���e�w� ����6��)��� =�_��F�X�j�|�K� ������������� 0BTfx�?�?�? ����3�,> bt����O ��//(/:/�� ��/��/��/�/�/  ?��/6?H?Z?l?�/ �?#?�?�?�?�?�?K/ ]/o/O�?hO�/�O�O �O�O�O�?�O
__._ QOR_�Ov_�_�_�_�_ OO1OCOE_*oyONo `oro�o�oe_�o�o�o �oo�o�o8J\n ��_�_�_o�;o �"�4�F�X�'|��� ����ď�i����� 0�B�����ɏ�� �ҟ������>� P�b�t�����+���ί������T_ER�R T���"�P�DUSIZ  j��^ɐ�9�>R�?WRD ?�Ō���  guest���������ȿڿ쿣�SCD_�GROUP 2UV�� ����1���!��2�ǒ  ,�C�	$SVMTR__ID 2�Ti�$GRP_2��$AXIS_NU�M Y�z�f�N�F��SV_PAR�AMiɑ� ,�$MOT_S��T�TP_AUTH �1V1� <!iPendan����Jũ���!K?AREL:*���KC3�C�U�+��VISION �SET��ߊ���! �߸���(������e�<�N��r����C�TRL W1���谡
��FF�F9E3�F�RS:DEFAU�LT�FAN�UC Web S_erver�
�� z����������������� �WR_CON�FIG X!��m��"�ID�L_CPU_PC�0���BȊ�K  ;BH1MIN<)�OGNh�O+�`����7�3 NP��IM_�DO��TPM�ODNTOL� >�_PRTY�K��OLNK 1Y1���#5GY�k}�MASTE� ���	OSLAVE Z1�����O_CFG��U�O����CYCL�E��*�_ASG� 1[l�
  ]/o/�/�/�/�/�/ �/�/�/?#?5?G?��0"��`�5�_��I�PCH/���RTRY_CN0����SCRN_UPD_��9� ����\1�&�O&��$�J23_DSP_�ENB�01�%�@OBPROC%C���JOG�1]1��8��d8�#?�R;�OR??U�S��LQ�O�O_#_�OG_Y_k_}_��'ҟ_[C�POSREEO�K_ANJI_�K�H�S1��3^���U<�_�UCL_L[ m2��?�PEYLOGG+IN�&��}A9���$LANGU�AGE m��e*� �a"�LG�2X��������x&Х��P���Q ���'�0������M�C:\RSCH\�00\�}`N_D?ISP `1���p���O�O �LOC��BDzj�A�cO�GBOOK a;+~@����q�q�pXCy������*�=�0�O���	 �u�y��Fu����!ua@BUFF 1b ��2��ڏ�r�� �����$�Q�H�Z��� ~�������Ɵ������ �M�D�V�����D�CS d�} =���L�����!������!���IO 1e;+ 
OZ����Z�j�|�������Ŀ ֿ�����2�B�T� f�zϊϜϮ����������
�5�Ez TM  2{d�_c�u߇� �߽߫��������� )�;�M�_�q����p����qw8�SEV�0�2}4�TYP@��R�3�E�W���QRS�? Ko���2FL 1fC��0�˯�������%7h�TP�_`@�"�k}NG�NAM%D�e���UPS*pGI�5a�5}�_LOADB@�G %2z%M�ANUTENTIONPINCE��D�$MAXUALRMm7�{8�'_PR�4�0�sM�C-pg;)[�q�s�Pc@P 2h�V ��	"���0���t�� ��� /ɨ/O/:/ s/V/h/�/�/�/�/�/ ?�/'??K?.?@?�? l?�?�?�?�?�?�?�? #OOOYODO}OhO�O �O�O�O�O�O�O�O1_ _U_@_y_�_n_�_�_ �_�_�_	o�_-ooQo coFo�oro�o�o�o�o �o�o);_J �fx��������7�"�[�D_LDXDISA� �B�3�MEMO_A�P� E ?��
 �c���ɏۏ�����#�5�IS�C 1i�� � M����b����L�՟�����J�C_MST�R j���SC/D 1k����g� 韋�v�����ӯ��Я 	���-��Q�<�u�`� ������Ͽ���޿� �;�&�8�q�\ϕπ� �Ϥ����������7� "�[�F��jߣߎߠ� ��������!��E�0� U�{�f�������� ������A�,�e�P� ��t��������������+O:s	�MKCFG l'��n�LTARM_*�m���q���,METP�U9d��/�ND�CMNTd�% � n'�c���{�%POSC�F1<PRPM�0�STOL 1�o'� 4@C�<#�
�n�/' �//1/s/U/g/�/ �/�/�/�/�/?�/	?�K?-???�?k1%SI�NG_CHK  y�t�ODAQ��p�=���5DEV� 	'�	MC}:�<HSIZE���C�Ȼ5TASK �%'�%$123456789 \O�nE�7TRIG 1	q`��%H��OA��O0�O�O)�>FYP)A�E��4�3EM_IN�F 1r�� `)AT?&FV0E0�Og]�)OQE0V1&�A3&B1&D2�&S0&C1S0}=V])ATZg_�_�TH�_�_vQ�Oo�XAo?o�_coJo�o�o M_�oq_�_�_�_ �_<so`r%o� Q�����o�o&� �o�o�on�y3��� ȏ�������"�	�F� X��|�/�A�S�e�֟ ����1��0��T�� x���q���a�s�䯗� ����,�>��b����� A�K���w��ǿ�� ɯ:�����#���G� ������ϡ����#��H�/�l��?NITO�RLG ?K  � 	EXEC�1j��2��3��4���5��@��7��8
��9j��6��� ������������ �����������2!�2-�29�2�E�2Q�2]�2i�2�u�2��2��3!�3�-�3�һ1R_GRP_SV 1s<[� (s1@����L=��->k�׮]�S��=�FA_D�,N�PL�_NAME !�S���!De�fault Pe�rsonalit�y (from �FD) �RR2�3� 1t)4�x�)4�����0@ dp*<N `r������ �&8J\n�82�������@�
//./@/�2<� j/|/�/�/�/�/�/�/��/??0?B?  � �\  ��  ��`��  A�  Bm0UTm0��0
Y0�]0~����  ��i0�h0Bm0pm0� � C�0C�0P �D�  D��N�2E@�2�2z�0 �1�0�1�2�0�9�2�0��6�4EK  E+� E��6�2�00�2 A DJZ��3A @DI�2�5�4�9�:�1;�7�:�5�@�5�O�;P�O�3�1�1E�1��0?�` E���G�4E���C�@Q�A@] Y$UP�5#V��D QL]hT�FQ8@�B U A U�T�R YU Q|UU�@�Y�Q�]�Q�Y �@B�YAP�1�R4o Bg�UXo�S�1Q`ong �Q�o�o�o�W�o�o�o� 2DV`tU0�DJxE�P/E�R�q�S2O��  l0��{q�d �sU0��}���tp�I<Z*����y�����`q�0 mb�T� @�5?h0p�T�?q�p�q�@u��5o����;�	l��	 � ���pXJ�����X � �? �, �ނO��K��K�z�K�ɜK@0>�KH�K$�@���������5��N��?��P�@'��6\����"��I�ڿ�
��}�v������X������0�/
=Âp¬0����  >ڃ��w�#�^���l� Y"�0��q����͔��,'��h���𗐿�  �T��  �`��v��	'� � ���I� �  ��-`�:�È~��È=���إ$�@���Z����Z��t'�5�o�yN��j�  '���O�?��@�t�@��@����X����Bd0Cf�0�pB��1��q��C�%
��e �_  ��^�/�B-`���$Ń�P���A�q��1ș_����oϕπϹ� �
��`��n� #�x�ݱ�� ؀���:m��q���?��ff��0��� ��d�v�%���.��?Y����|��	(q���P�����ȃ�Ȅ2�?33��������;��;����;�D�;��$;�< J!l �=�L�~�Z����=�?fff?��?y&zࡔA���@�,��j��u� ����p���n���^約 O�$��H�3�l�W����{���������+���F-���&��J��k���=�ɘD�@�|���0�  F�� ����5 Y DV�z�ƚG�� �/a'/�N/�r/Є/�/�/G�A�0����O�tp��B�0h/?�d/%??I?4?��-�A �0t2-`|1�?�u�?\?�2;囏Ŝ?�ؠ�?�?OO*�į���W*OC��@�` #Ca'O*�4��0�1��A��ܨ���C�>CR BA�Aˉ7�����"���z���q���=�\)xO� ʊ�=��=qA�B){���O~� �(��g�/P��qBp��߿{��8R��K���J?&DK���	HwW�H�'��!��LA��L�9K���4HŀHH�� h_zP��L�m�J�sdHK�� H-�A� �_wO�_�_o�_%oo Io4omoXojo�o�o�o �o�o�o�oE0 iT�x���� ���/��S�>�w� b�������я������ ��=�(�:�s�^��� ������ߟʟ�� � 9�$�]�H���l�����ࢯۯƯ���G�$�� C���4�F@�؇�u�8�V��0��������Ͽп�����?��F( Q�g`��G� ���xŎ8E�Y��>x�	3�Z�_�Ϧϴª�����ϰ�fC3�g���̅����3�Ȭ ��X�F�|�jߠߎ�J�5P��P�������N�����.����P�b����7(���C@�C@5��� �
�@�.�d�����`������������0������&�  JK  � @^��v������2 D�J�E-���0��B}1q1�}0C�f@�AC@@��?FC@J�m��C�B���z���3��wE�(��F����
//**@9$��J�4C@C@���4�;
 */�/�/�/ �/�/�/�/??/?A?`S?e?w?�J�2��������$MS�KCFMAP  �D� �g!c!�>�3ON�REL  s���1�а2EXCFENB�7
�3�5A�FNCODJOG_OVLIM�7d@�Bd�2KEY�7�eE�2RUNUL�eE�2SFSPD�TY��FE�3SI�GN�?DT1MO�TWOA�2_CE_GRP 1zD�3\,�;_$�__ q_�[_�_S_�_w_�_ �_�_o�_oPooto �o=o�oao�o�o�o �o�o:�o^pW��K������1Q?Z_EDIT�D�7��3TCOM_CF/G 1{�=r&I��[�m�
)�_ARC�_B��DIUAP�_CPL��(DNO�CHECK ?�; ����� ��
��.�@�R�d�v� ��������П����;�NO_WAIT_�L�G�	PNT1��|�;i+F�_ER�RQ2}�9�ф A�����ï���3x���ńT_MOt�}~{�x G�V�|D��8�?\�_�I�b 6�m�PAR�AMu��;��f&4���w� =�� 345678901'�9�K�"�j�|� Xψϲ��Ϡ��������w�,�>�ѿb�ƃ�UM_RSPAC�E�?R�o��ߥ��$?ODRDSP���F�$HOFFSET_�CAR�����DI�S����PEN_FILE��Ao�����PTION_IO�vO�A;�M_PRGw %��%$*t�����WORK 5�W'C ���D�6��2���S���	 �a���6�C����RG_DS�BL  DC�j,@���RIENTTO�0���2 ���UT_SIM_EDC��2�2��V��?LCT �P�����ݒ�_PEXE���RAT��\F$E�����UP ���x E �/A'�es	�$��2St�)4�x)4��>��@ dRߺ ���&8J \n������ ��/"/a�2�R/ d/v/�/�/�/�/�/�/�/��<A/?0?B?T? f?x?�?�?�?�?�?�?��?�����)P� � ��  �p�A��  B!@�B��Y@H@��  ��@p�BJ!@p!@�d�c����P D�  D;��bBE@jB_Bzd�`A`@{A{Bx@�I�{Bd@�F|DEK  E+� E��F��Bx@kB�A�D�JZ� fC�A�D�I�B�ElD�I�JlA;eGJ�E<P�E@c_}Ks_aC[A{AEhA��m@�` E��\�WxDE���S��@ �Q�Q�]�Y�U�P�E�V��T�Q md�V�Q�@ �R�U�A�U@dcb�Y�U�Q0e�U˵@�ida�m da\i<P�B�i�A�P[A �b�o�g�e�chA�Q "wda4Bp�gx ������
����"� @E�W���P�s���j�����(�(��� O 1y(ӿH(�&���`�0�� @�Eo�o���?|�C@�E��.� _ ;�	lo�	��� ����pX̰��q���X � � ��, �����H���H��H��PuHV�2H�H_3��<������B�!@	�C`���@�γ�4@�L@�
=�g���`@D�(�:�L�)�A�ߟ�½��ªVy�H@����p�ˣXQ�ϡ�hD��D���  �  ������Q�6��%�	'� � �T�I� � � ��`R�=��q�x���(�@��@�����ʿ;��$��߯�'�Np�"�  Q'F�:ą�Ca�B@Cfd�B�Au�G�Y�� ��  ��C�%  �*��^��/V�B�`��8p���;� ���� ��wA���^�'�M�8ߜqߨ�
�`��U�?n� �x����2�� ����:O���}Q��?�ffǏ�����z߶�%�ㅡ8���E�S�?Y����$4�|�(����P����ő������?333�Q����;��;����;�D�;��$;�<� Jl�����6��޳8���?fff?淰?&2�A�=D�@�,P�Q� ��-�9�T�(���&��� �l������ ��$ H3l~i�� ����s������,V��Dڹ@�U�@�  Fg�D� �����/�/ G/2/k/�����-]/�/ �/=?y/*?<?N?4`?��AL@��j��	�d�B8@ ?�??�?`�?O�?B�'�A�*D �`4A;O�0�?bO����<S�}�?�؏O�Oh�O�OQ��g��W�O�C��P�` Ca��O�*�D��@�ALQ@�I	�b���C�>CR BA�Aˉ7���Q��"���z���q���=�\)0_�0ʊ�=��=qA��B){�녨_~�0�(��g��P��qBp��߿{��8R�MK���J?&DK���	HwW�H�'��1�MLA��L�9K���4HŀHH��  o2`��L�m�J�sdHK�� H-�A� Jo/_�o�o�o�o�o�o �o%"[F j������� !��E�0�i�T���x� ��Ï���ҏ���/� �?�e�P���t����� џ�������+��O� :�s�^�������ͯ�� �ܯ� �9�$�]�H��Z���~����KG�$��ſ C�����@��?�-��V��07�>�w�b���ψϠr��Ͼ��ϲV(xA�g`���ϸ���0Վ�ųY«N0߲S3�Z�_L�^�lҪ��xߊ߰�fC3�g�߶܅����3�Ȭ �������4�"�X�F�J�EP��P��!�/���߿������`�����S�>�V�7(`�r�{�{5��V� ������������/`I ��JXj�t0���������  JK  � �@.dR�r��2 D��E-��0�VB5A)A�5@C�P��A��@`9O�/"/2,C�����2/[/i*�CN�E;�(�VF�i/�/H�/�/�*@�$�XxD%����O�|D�K
 �/E?W?i?{? �?�?�?�?�?�?�?O�O/O�ZB��\�����$PAR�AM_MENU �?���  DE�FPULSE;K�	WAITTMO{UT�KRCV�O� SHELL�_WRK.$CU�R_STYL�@��LOPT��OP�TB�O�BC�OR_DECSN�@{�N\ H_Z_l_�_�_�_�_�_ �_�_�_%o o2oDomo�hASSREL_I�D  +�x�@}dU�SE_PROG �%wJ%io�o}cC�CR�@+�C�g_HOST !wJ#!�d#�jT���o�?sqAs{�k_�TIME�B�f�e~h@GDEBUG�`�wK}cGINP_F�LMS�~�xTR\��wPGA � �|�N��CH��xTWYPEtL� ho bo������Ώ��	�� �(�Q�L�^�p����� �����ܟ� �)�$� 6�H�q�l�~������� Ưد���� �I��uWORD ?	&��	RS���PNS��D��J9OQ�TEbpF��TRACECTL� 1���A� ��% &e��� ߾��DT �Q���ӰD� � 
 ��������Ď`!��*��	�
�Ϡ0�B�T�f�x�z���� y�0y�0y� 6�y�0y�0�ϻ�����C���C���:� L�^�p߂ߔߦ߸��� ���� ��$���;�-� _�q��������� ���S�%��)�[�m����ã��£��� ��ң�ң�ң�� ��&ң�£��£��� ��~£��£��£�� ��£��������	 -?Qcu�� ���������� ߺ��φϘϊ�� �����S_/q/ �/�/�/�/�/�/�/? ?%?7?I?[?m??�? �?�?�?�?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_�_�_�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]o� �������� #�5�G�Y�k�}���[/ ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�W� i�{������������� ��/ASew ������� +=Oas�� �����//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?#?5?G? Y?k?}?�?�?�?�?�? �?�?OO1OCOUOgO yO�O�O�O�O�O�O�O�	_Q�$PGTR�ACELEN  �Q  ���P�'V_U�P ����2VQ^PBQWP'Q_CFG �VUS@SQWP��T�9P�_�\kRDEF�SPD �v\lQ9P�'PINnP�TRL �v]�P8�U�QPE_C�ONFIrP�VUO�VQ�T�Y.'PLIDoS�v]�Q~EaGRP 1�g����QC%�  �ᙚQA��=qGY� G�cX Fg@ A��  D	��T	�Pd�T�i�i5a5`?� 	 �_�R�[�o ´s�o�kBp>qT>�x�rH9B!ၖ��~� <T?��<]/�� ��U�@�y�d����@����я��⏠`z�%�P
�M���]��� n�����˟���ڟ� ���I�4�m�X������!Q
V7.1�0beta1�V� @�p�@z?=q@��R�aʡ�C  C5PB|�ܣDf@ �C���`� D�� D� C�`f�`B�䠃`C/�`p�R�r�`1�C�U��$�BdKNOW_M�  �U~VBdSV� �mi�-e:�ſ׿�z��@��
�CσR�mAcMfc)���8Plڢ	�Rܡ�  �b�� ^ ����S��ˠ`���IˮiRLMRfc�y�T�z��QCz����u�8�J�6mSTfa1 {1�V[
 0-e��$բ�  �ߙ߫� ��������4��)�;� M��q��������@�����T�h�2s�9��Q�<��a�A3r�������l�4��������l�5"4Fl�6_q��l�A7����l�8�p!3l�MAD3V� ^Vh�PARN_UM  V[2�\�j�SCH� ^U�
�� )@S%UP�D���e\/�_C�MP_o�3PWPP'�WjS_ER_CHK�%|X�&/�+�RS�}�Ba_MOȜ�/�%_�/\e_R�ES_GrВv�  ��nr?e?�?�?�?�? �?�?�?OO8O+O\O OO�_44q�><N?�O 35��O�O�O53 �O �O _53^ _:_?_53 � Z_y_~_53� �_�_��_53K�_�_�_52V� 1�v�$1��@�c���"THR_�INR0"!W�(5d�kfMASSxo Z�gMNwo�cMON�_QUEUE ��v�	6#0/��TN�y U�!N�f�+�`E�ND�a?yEXE(u> BE'p	�cOPTIOw&;�`�PROGRAM %�j%�`6o�~�bTASK_I��o~OCFG ���o���DATA�rÖ�@0�2 ��t���������g��� ���(�ӏL�^�p����5�INFOr×Q���d=�ڟ���� "�4�F�X�j�|����� ��į֯�����0�hB������Q� lI��� DIT �����5�WERFL�Ix^ci�RGADJ� ���A�  b��?#0�d�RG�a���y��?9���a�<@���ɖ�%ah�ϸ���2�����`\hF�]b2�2�A(d�t$���*��/�� **:��#0����v���������W�Ab5�Ac	��-� ?߬�c�u߇ߙ��߽� ����N�I��)�;�� _�q���������� ����%�7�I�[�m� ��������������� !�EWi{� ����/� ��Sew��� ����//+/U/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]?�? 	 ��?�?O�7 ��9O��OfOO�O�����PREF ��%�OpOp
۵IOORITY�g��߱MPDSP�qͿ�G�U�g��ڶOG��_�TGʰ�r�j*RTO�E�`1��� (/!AFs`E�`s_~~W!tcp~_>�]!ud�_�^?!icm�_8o�+QXYà���Oq)� ��2oDoOp�,omoPe\o�o�o �o�o�o�o�o�o;@M4qX��*)S�â�MU�����?W!�}�6��/�Ɉ�K�V��~ȁƺ�A~G�,  ��@ w�������͏�E�t�CᣴO�Cղ߱POR_T_NUMS�����߱_CAR�TREP�@����SoKSTAW J�SAVE ���	2600H738҈O�Or�`������LÉ7�����7Z�URGE_�ENBʹ��aWFF(�DOV{�EVWlP�I�ձ)�WRUP_�DELAY ����=�R_HOT �%�ֲ=�ɯZ�R_NORMAL���򲸯�ܧSEMI���Q���QSKIuPȓ��� x}O ��yO��̿޿���=� ����4�F�X��|�j� �ϲ����Ϝ������ 0�B��R�T�fߜ߮� �߆��������,�>� �b�P����p���������(�2��$�RBTIF7_�AR�CVTM[BT��E�DCRm��t�� Э�E8����Ed��C���B��\8������P(GŃ�#��Añ��\7�´B������ ;���;���;�D��;�$;�< Jl��Se ������� ��	-?Q�G�RDIO_TYP�E  ϝG]E�FPOS1 1���
 x?��Z@ �</�^��/v/ a/�/5/�/Y/�/}/�/ ?�/<?�/`?�/�?? 1?C?}?�?�?O�?&O �?JO�?GO�OO�O?O �OcO�O�O�O�O�OF_ 1_j__�_)_�_M_�_ �_�_o�_0o�_To�^�2 1�����oJo�oFo�ojo�3 1��o�o�o�o`�K�S4 1� +=w����S5 1��������u���,�S6 1�C�U�g����
�|C���S7 1�؏����6�����؟V�S8 1�m����˟�I�4�m��SMAS/K 1�z ��������XNOw��x����MOTEL��۫��_CFG ���b����PL_RANG�O�Q�OWER �����#�SM_DRYPRG %��%�����TART� �|�ʺUME_PRO����&���_EXEC_EN���ĄW�GSP�D��A�Iȓ�X�TD�Bd�v�RM��v�MKT_��Tw��E��OBOT_ISO�LCخF�2�b����NAME ��ÉOB_O�RD_NUM ?�|��H�738 ~  ����r���}�y� �2�Dr��h�z��r� �����r����
�r��x+��PC�_TIMEg�S�x�E�S2320�1������LTEA�CH PENDA�Ni�,���7����PMaint�enance C�ons��$�"���TKCL/C�ٰp����o� �No Use��N��9���NPO���^���Y����CH_L������	=��MA�VAILSѸ�K������SPACE1w 2�� �@K�����2���K�L��b���8�?� ����IjA z���������' :�_pW�� �����S' /:/�_p/W/�/� ����//#/?6? �/K?l?S?�?�/�/�/ �/�/�??1?3?�?GO hO?OQO�?�?�?�?�? �OO-O_}OC_d_v_ ]_�O�O�O�O�O�__ )_o<o�_a_roYo�o �_�_�_�_�oo%o 8�oMnU��o�o �o�o�o�o�z� I�j�A������ ����/�!��E�f�Px�O�a���2���� ��͏ߏ���%�4�U�@�j���r�����3�� Ɵ؟����� �B�Q��r�5�����������4 ѯ�����ǿ=�_� nϏ�RϤ��Ϭ��ϥ�5� ��$�6���Z� |ϋ߬�o�����������6��/�A�S�� wߙߨ�������������7(�:�L�^�p� ������������1��8E�W�i�{� ��;�������9 N��G �Ne E�
�7 �  e� ��//%/7/g��V-�c�/+�/�d � ���/??&?8? J?\?R/d/v.g:�?�; �?�/�/^?O*O<ONO `OrOh?z?�?�?�?�O �O�?�?~O8_J_\_n_ �_�_�O�O�O�O�O�_w `F @� �+e�/9o_Ywa�U o�o�o�_zj{o�o�o �oI[%/ As�w���� !�?��'�i�{�E�O� a���Տ���\
Yo*����_MODE  ye@�S �e��_�Z�Uo~��П��	�� �CW�ORK_ADP�
�^dȡR  �er g��Q�_I�NTVALP����[�R_OPTIO�N�� [��V�_DATA_GR�P 2��XpDPP������ C�1�g�U���y����� ����ӿ	���-��Q� ?�u�cυϫϙ��Ͻ� ������'�)�;�q� _ߕ߃߹ߧ������� ��7�%�[�I��m� ������������!� �E�3�U�{�i����� ������������A /eS�w������W��$SA�F_DO_PUL�S;�X��AZ�1!C?AN_TIMO�!U���BR �(��C�(�f0�"�����Ē����S ���� �//�7/I/[/m/X/�/���C,"2�$��d�(�!�!�&�@�\
??�.?*��)�/ ߠC4��_ 3b  �Tf�W?�?�?�?�9T D���?�? O O$O6OHOZOlO~O�O �O�O�O�O�O�O_��<���%_X_�j_'Y+a��Q;��o*���p(]
�t� �Di���� -��,"���Q ��y�_o o2oDo Vohozo�o�o�o�o�o �o�o
.@Rd v������� ��*�<�N�`�r��� ������̏-��T?�� ��+�=�O�a�s��� ԏ�%��ß՟������/�A�S�X���-�0 R2�S�U�]����ȯگ ����"�4�F�X�j� |�������Ŀֿ��� ��0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�t�ߏ�ߪ� ����������(�:� ��^�p������� ����Y�����,".�@� R�d�v����������� ����	'9K] o������� �#5GYk} ��������X�$_�3/C/U/g/y/ �/�/�/�/�/�/�/	?@?-???Q?c?q:0/�z?�?�6������?�=	1234�5678�R !�B�P
�8.  �PO)O;OMO_OqO�O �O�O�A//�O�O�O_ _*_<_N_`_r_�_�_ �_�_�_�_�_m�O$o 6oHoZolo~o�o�o�o �o�o�o�o 2DoBHU}�� �������1��C�U�g�y�����k;�j��ӏ���	� �-�?�Q�c�u����������ϟ��
iD� ��%�7�I�[�m���� ����ǯٯ����!� 3�E�oi�{������� ÿտ�����/�A� S�e�wωϛ�Z����� ������+�=�O�a� s߅ߗߩ߻������� ���'�9�K�]�o�� �������������#�5�G�$@d�v��[�������)"C�z  A�*   �(2�4A���A!��0Ě22�b�I[m���0/���8�� �!3EWi{ �������/ ///�S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�?��$SCR_GR�P 1�(ӈ��(ӑ ~@t ��
 �1 	 �3  AB	D��"M�7GpJO8OqO��� ~nBD�` D���C�GnK�R-�2000iB/1�65F 5678�90. �DX. �R2D7 �@B#
1234�EAFnAZ� CV�1�B&�3�1�nAJBATY	ER�_�_�_��_�_�\��H��0�TG�2&o5O@6o\ono=FM/
Io@�oEo�o���o��h,P��TpE  p��AB���B��ffB�33B�K  +v�5wAA���G  @
 _uA@<�@o  ?��wr�H-p�JzAF@� F�`�r�=GC�  ��� �� D�/�h�S���w�7q_q��r������ʏ܄B� ��0��T�?�x�c� u�����ҟ��������*��CZOH�m����  j���
�q@�r�AO��=G��߯-p���W\NCa�5�B$AA�G�1Z��o�e �Y�
 {������º��׸���Ŀ P�(!�'�9�K���1EL_DEFA�ULT  XT�_�
 _��MIPOWERFOL  ��w���gWFD n� w��^�RVENT 1O���`u����L!DUM_E�IPM����j!?AF_INEk�ߞB$!FT��>���b�!"o�� ��Q߮�!RPC_OMAIN�ߖ��ߜ����VIS�ߕ	����F�!TP9�P�U=���d5��!
�PMON_PROXY����e����Y�����f��*�!R?DM_SRV+���9g�v�!R!T�����he���!
��M�����i��!R�LSYNC5	�8��Z!ROS��ρ�4I�!
�CE[�MTCOMd���k��!	�OCONS���l� >u�b9�/A�� w����/�@/�//+/�/O/a/Q�R�VICE_KL �?%�� (%SVCPRG1�/D:�%2??� 3+?D0?� 4S?X?� 5{?D�?� 6�?�?� 7�? �?� TO<9O K�$��HO�!�/pO�! ?�O�!E?�O�!m?�O �!�?_�!�?8_�!�? `_�!O�_�!5O�_1 ^O�_1�O o1�O(o 1�OPo1�Oxo1&_ �o1N_�o1v_�o1 �_1�_@B1�_�/ �"� �/� ��1� ����@�+�d�O� �����������͏� �*��<�`�K���o� ����̟�����&� �J�5�n�Y���}��� ȯ���ׯ���4�� X�j�U���y�����ֿ ������0��Tϖz_DEV �ɿ�MC:\� w
�n�OUT`��h��j�REC �1ŭuh��� �� 	 \�������3�lu:��c��n�
 �Tpvj�6 sS�� � ����  _�  Пл�u\��X�r 1��h�e=h���ů� ���U�h�+h���2���������'�M�;� q�_��������� ����#�I�7�m�O� a������������� !E3UWi� ������ A/QwY��� ����/+//O/ =/s/a/�/�/�/�/�/ �/�/�/'??K?9?o? �?c?�?�?�?�?�?�? �?#O���O)OOQO �OuO�O�O�O�O�O_ �O)__9_;_M_�_e_ �_�_�_�_�_o�_%o 7oo[oIoomo�o�o �o�o�o�o�o3! WE{�o��� ����/�A�#�e� S���w��������ŏ ����=�+�a�O��� ��y�����ߟ͟�� �9��I�K�]�����෯��ۯ�׽�V 1���� (ӯ&���TOP10 1���
 ��,�v������@�YPE��l�H�ELL_CFG ��{�h�	� � ��B�RSR��/�h�Sό�w� �ϛ��Ͽ���
���.���R�=�v߈ߚ��
����%�����ߨ����������S��װ�2h�d��|��϶HK 1�ݻ 
����� ����������+�=� f�a�s������������h�϶OMM ��ݿβFTOV_�ENB���ƺOW_REG_UI=~ͲIMWAIT:���mOUT^��o	TIM^����VAL~p_�UNIT9�ƹL]CW TRY^Ƶ���MON_AL�IAS ?e	�he�Vhz� ���R���/� %/7/I/[/m//�/�/ �/�/�/�/�/?!?3? E?�/i?{?�?�?J?�? �?�?�?O�?/OAOSO eOwO"O�O�O�O�O�O �O__+_=_O_�Os_ �_�_�_T_�_�_�_o o�_9oKo]ooo�o,o �o�o�o�o�o�o# 5G�oX}��� ^������C� U�g�y���6�����ӏ ������-�?�Q��� u���������h��� ��)�ԟM�_�q��� ��@���˯ݯﯚ� � %�7�I�[������� ��ǿr�����!�3� ޿W�i�{ύϟ�J��� �����Ϥ��/�A�S� e�߉ߛ߭߿���|� ����+�=���a�s� ���B��������� ��'�9�K�]�o���� ������������# 5G��k}��L �����1C�Ugy#�$SM�ON_DEFPR�O ����� �*SYSTEM*�  ȏRECA�LL ?}� �( �})cop�y mdb:*.�* virt:\�tmpback\�=>portuc:14768 &`/&/8/J/#}/��frs:orde�rfil.dat��emp�753�2 /�/�/�/Z$'b&*.dv/�'�/?�-???R,
xyzrate 61 �/@�/?�?�?�?Y%b7��,{?�?O0OBOU)0��:manute�ntion.tp�o?�&O�O�O�O[#2 b/t(�B_&_8_J_ ]!��OD_�_�_�_6T*-x�D:\k_�P@�,�_!o3oEoX&.�Ua�_�_2 o�o�o �o�O�Ot_�_ 2D W_i_{_���U/��ozO:18700 �#�5�G��/�/� 
�������R?d?v��� �+�=��?�?���� ����UOgO������ $�6�H��o������ ����ʯ]x����� /�A��_�_yo����� ��ſXojo{�����"� 4�F�Y�k�����ϲ� ��ׯ������0�B� U�g������߮���ӿ �v�	��,�>�Q�c� uχϘ���O���|� ��(�:�L�_��߃� ����������n���$6H[�1k���О���y9�np�inceauto ����!3EXj�� ���Ugy� /./@/ӟ� /�N/ �/�/�c/�~/�/*? <?�/a�??�?�? �?�q?�?�?&O8OJO ]?�?OO�O�O�O[� m���O&_8_J_���O�/_�_�_�_�"��$SNPX_AS�G 1������Q� P� 0 '%�R[1]@1.1,�_i?��#%oDo 'ohoKo]o�o�o�o�o �o�o�o�o.8d G�k}���� ����N�1�X��� g�������ޏ���� ��8��-�n�Q�x��� ��ȟ��������4� �X�;�M���q���į ���˯ݯ��(�T� 7�x�[�m�������� ǿ����>�!�H�t� WϘ�{ύ��ϱ���� ��(���^�A�hߔ� w߸ߛ߭�������$� �H�+�=�~�a��� �����������D� '�h�K�]��������� ��������.8d G�k}���� ��N1X� g������/ �8//-/n/Q/x/�/ �/�/�/�/�/�/?4? ?X?;?M?�?q?�?�? �?�?�?�?OO(OTO 7OxO[OmO�O�O�O�O��D�TPARAM ���U�Q W�	��JPXTXP��XOFT_KB_CFG  %S��U?TPIN_SI/M  �[4V�_�_�_7P�PRVQS�TP_DSBn^�4R�_"X�@SR ��qY � & ��_/o%P<VTH�I_CHANGEw  %T\W~OaGRPNUMOV� djOP_ON�_ERRYhZY�aP�TN qUc`�AKbRINOG_PRy`�n�@wVDTsa 1�Ya`  	8W"X 0BTfx�� �������,� >�P�b�t��������� Ώ�����(�:�a� ^�p���������ʟܟ � �'�$�6�H�Z�l� ~�������Ư���� � �2�D�V�h�z��� ����¿Կ���
�� .�@�R�y�vψϚϬ� ����������?�<� N�`�r߄ߖߨߺ��� �����&�8�J�\� n������������ ���"�4�F�X�j��� �������������� 0WTfx�� �����, >Pbt�������?SVPRG_�COUNTOV�8�a^U"ENB�o	%�M3#|eA/UPD �1�kT  
 �%R�/�/�/�/�/�/ �/??,?>?g?b?t? �?�?�?�?�?�?�?O O?O:OLO^O�O�O�O �O�O�O�O�O__$_ 6___Z_l_~_�_�_�_ �_�_�_�_o7o2oDo Voozo�o�o�o�o�o �o
.WRd v������� �/�*�<�N�w�r��� ������̏ޏ��� &�O�J�\�n������� ��ߟڟ���'�"�4�� +YSDEBUG� y �J�da)l�S�P_PASS%�B?~�LOG ��x%c#J��G�T�  �]!J�
MC:\��Z���_MPC��x%,�>��x!�\� x!�S_AV ѳ�Фl�J��SV_��TEM_TIMEW 1�x)��(Ѡ�áСȯ)T1S�VGUNSs %'�a%�	�ASK_?OPTION x%t]!'!)�_DI���4/E�BCCFG 3�л�� ������`��������� �����7�"�[�F�� jߣߵߠ��������� !��E�0�B�{�f�� �����������J�	�8�
�k�}���Z� ����������c�;� ��#I7m[� ������3 !WE{i��� ����//-/// A/w/](H��/�/�/�/ �/]/?�/?9?'?]? o?�?O?�?�?�?�?�? �?�?�?OGO5OkOYO �O}O�O�O�O�O�O_ �O1__U_C_e_g_y_ �_�_�_�/�_�_o-o ?o�_coQoso�o�o�o �o�o�o�o)M ;]_q���� ����#�I�7�m� [��������ŏǏُ ���3��_K�]�{��� ���ß��ӟ���� /�A��e�S���w��� ������ѯ���+�� O�=�s�a�������Ϳ ���߿��%�'�9� o�]ϓ�I��Ͻ����� ��}�#��3�Y�G�}� �ߡ�o��߳������ ����1�g�U��y� ���������	���-� �Q�?�u�c������� ��������;M _���q���� ��%I7m [}����� /�3/!/C/i/W/�/ {/�/�/�/�/�/�/�/ /??S?	k?}?�?�? �?=?�?�?�?OO=O OOaO/O�OsO�O�O�O �O�O�O�O'__K_9_ o_]_�_�_�_�_�_�_ �_o�_5o#oEoGoYo �o}o�oi?�o�o�o �oC1Syg���v�p�$TBCS�G_GRP 2���u� � �q 
 ?�  ����� @�*�<�v�`������r��s��|d0�ہ?�q	 HDw)̪�&ff�����B\�r�!��'333?���!�#��L�͇�L������C�����ϖ��CA�C4 ����Ř@�� ����HŘ���HA���@�p ������¯�����
��կ�5�R�a�7�p � ,	V3.�00�r	r2d7a�	*�����rЬ�k���(�p7� �㰵��  ������M�&�-ÿqJC�FG هuX�q�-��W���9-ς���Ϩ� �ʐp������ ���$� �H�3�l�W�iߢߍ� �߱���������D� /�h�S��w����� ����
���.��R�d� �r�`o�����=����� ������ D/h z��Y���� ��q�A�QS e������/ �/=/+/a/O/�/s/ �/�/�/�/�/?�/'? ?K?9?o?]??�?�? �?�?�?�?�oO)O�? IOkOYO�O}O�O�O�O �O�O__1_�OA_C_ U_�_y_�_�_�_�_�_ 	o�_-oo=o?oQo�o uo�o�o�o�o�o�o )M;q_�� �������7� %�[�I�k���;O���� ͏w������!�W� E�{�i�����ß՟�� �����-�S�e�w� 1�������ѯ����� ��)�+�=�s�a��� ������߿Ϳ��� 9�'�]�Kρ�oϑϓ� ����������#�5�ߏ M�_��ߡߏ��߳� ���������C�U�g� %�w���������� 	����?�-�c�Q�s� �������������� )_M�q� �����% I7m[}�� A���/�3/!/C/ i/W/�/{/�/�/�/�/ �/?�//??S?A?c? �?�?�?g?y?�?�?O �?+OOOO=O_O�OsO �O�O�O�O�O�O__ _K_9_o_]_�_�_�_ �_�_�_�_o�_5o#o Yoko/�o�o/Qo�o �o�o�o/UC y��[m��� ��-�?�Q��u�c� ������Ϗ����� �;�)�K�q�_����� ����ݟ˟���7� %�[�I��m������� ٯǯ��wo�o'�9�� �W�i�����ÿ��� տ��/�A���e�S� u�wωϿ������ϯ� ��=�+�a�O�q�s� �߻ߩ��������'� �7�]�K��o��� ���������#��G� 5�k�Y�����K����� ������1AC U�y������	�-Q;  9w{ {��{�$TBJOP_GRP 2�C��  �?�{	������K�� `p�p� ��?� � � {� @w�	 ߐD)�+%C2?
C랔{��G"333O!>����K/! LY p$<���d+!? !p$B`�  A�A$��� ��'+/=/O%O"�/�*�<+�~-C  B�{@!/?�/��/F'p%�%p=���5<ҙ*"P!p!��Cz!0�$�?�;C��6���C�p��.�?K�%p �;��:CA�4�"P$C�C4�?VO��?�?m(�Oj;(A�=)�/JhAH�0 YO�OpiO{O_+^fff?U<:f�/F !�0?B �@f_x_+_�_�Y�_�_ �_�_o�_�_!o;o%o 3oao�omo'o�o�o�o��o�o"�D�{�  ��G%	V3.0}0�r2d7��*mp�v{�w� GO �~d�� G�0G�� �G�| G�: �G�� G�� �G�t G�2 �G�� Gݮ �G�l G�* G�� HS�r�Fj` �~� �F�q � GX� G/� GG8� G^� Gv� G�ĺs�4 �G�� G�� �G�\ G� �=p =#�
|8�(1Cq�j�k�}�{��?�X���~�ESTPAR�p�o��HRրA�BLE 1ݵ$��{���� ��v�
������z���	��
�����{U�������'RDI����!� 3�E�W�i�єOٟ�@����+�=��Sן� �����"�4�F� X�j�|�������Ŀֿ �����0�B�TϚ ֠گ	���~������� `�r����������{¿NUM  CU� � ��̐�_CFG ��d��!@�IM?EBF_TT܁�8�逦�VERʓ��z����R 1ߵO 8x{v2� F��  �� %�7�I�[�m���� �����������!�3� E���i�{����������������_b̐/ �  k�Ԭ��T��6����9��I��/� �LTA_�b6���L�6���B���^�� 7��\��/ 
��:Q��);^���g]o  ��R�ƙs/ V�dà��/ Wش���
�/ [X�s%�H	/���_^���@���ӀMI_CHA�N�� �� �#DB/GLVL����ҁ�� ETHERADW ?��� ���������/?ˈ� R�OUT��!��!�54S?&<SNMA�SK�(���!255.�5Ys�?�?�?Ys�ӀOOLOFS_�DI�pM%�)OR�QCTRL �$�ɖ���1NT OUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_��\O�_�_�_ЃPE?_DETAI�(�:�PGL_CONF�IG �d�tф��/cell/�$CID$/grp1�_FoXojo|o�oD��?�o�o�o�o �o7I[m�  ������� �E�W�i�{�����.� ÏՏ�������A� S�e�w�����*�<�џ@�����+���}�� a�s���������)ѽ_�­����*�<�N� `�r���������̿޿ ���&�8�J�\�n� ��Ϥ϶��������� ��"�4�F�X�j�|�� �߲����������� 0�B�T�f�x���� �����������,�>� P�b�t�����'����� ������:L^ p��#����� $`�EU�ser View� 4oXjI�}12�34567890 �������@ ,c/��;2q=/ O/J�s/�/�/�/�/�/=�//C3�/!?3? b/W?i?{?�?�?�?�/�/<4�?OOF?;O MO_OqO�O�O�?�?<5�O�O�O*O_1_C_@U_g_y_�O�O<6�_ �_�__oo'o9oKo]o�_�_<7eo�o�o �_�o�o/Apo�o<8I���o������%�TF� ��ECameraFx������@��ҏ�����E�� 9�K����x������� ��ҟ�`�+/�'��� K�]�o��������ɯ ۯ�8��#�5�G�Y� k�2�pu`�?��ÿ� �����/�Aϸ�e� wω�Կ�Ͽ������� �~����?M�_ߞσ� �ߧ߹�����T��� %�p�I�[�m���� ߐ��O����:��1� C�U�g�y��ߝ����� �����	-?�� ���_������� ���9K]� ������R�� �o!/3/rW/i/{/�/ �/�/(�/�/�/D/? /?A?S?e?w?���� �?�??�?OO)O;O MO�/qO�O�O�?�O�O@�O�O__�?��9!_ Z_l_�O�_�_�_�_�_ �_aOo o2o}_Voho@zo�o�o�o'_qt	a�0�o�o	Ho-?Q cu��_��� ���)�;�M��o�l1Y������ɏۏ� ���#��G�Y�k��� ������şן�`��l2��/�A���e�w��� ������6�����R� +�=�O�a�s������l3��˿ݿ���%� 7�I�[�үϑϣ�� ���������!ߘ��l4-�g�y߸ϝ߯��� ������n��-�?�� c�u�����4��l5����T�9�K�]� o�����
������&� ��#5GY���l6e������� /��Sew� ������lz  w	+/=/O/ a/s/�/�/�/�/�/�/�+   /	/'? 9?K?]?o?�?�?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_ y_�_�_�_�_�_�_�_�	oo-o?oQoco�, � 
s (  �> ( 	 so�o �o�o�o�o�o% '9o]���}j: �K��  ��D�V�h�z����� u�ȏڏ�3��"� 4�F�X�j��������� ��֟�����0�w� T�f�x���������ү ���=�O�,�>�P��� t���������ο�� ��]�:�L�^�pς� ��ۿ������#� �� $�6�H�Zߡϳϐߢ� ����������� �2� y�V�h�z��ߞ���� ������?��.�@��� d�v����������� ��_�<N`r �������% &8J\��� ������/"/ i{X/j/|/��/�/ �/�/�/�/A/?0?B? �/f?x?�?�?�?�?? �?�?OO?,O>OPObOptO�O�?�p@ �B��O�O�O�C�G�`����O_&_8_J_\_ n_�_�_�_�_�_�_�] _o o2oDoVohozo �o�o�o�o�o�o�_
 .@Rdv�� �����o��*� <�N�`�r��������� ̏ޏ���&�8�J� \�n���������ȟڟ ����"�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ������I(A ��O�$TPGL_�OUTPUT ���1�1 ���,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p������������� � 2345678901����%�7� I�Q��2��x������� ����j���,>P��}Z���� �bt $6H Z�h����� p�/ /2/D/V/�  /�/�/�/�/�/�/~/ �/?.?@?R?d?�/r? �?�?�?�?�?z?�?O *O<ONO`OrO
O�O�O �O�O�O�O�O�O&_8_ J_\_n___�_�_�_ �_�_�_�_o4oFoXo jo|oo�o�o�o�o�o�o�o��}��0BTfx��}@�Ͽ�|����( 	 �� ��*��N�<�r�`� ������̏����ޏ� �8�&�H�n�\����� ����ڟȟ����4��"�X���OFF_�LIM#��������t�N_S]Vx�  �����P_MON ��َ��������ST�RTCHK ��Պ�-��VTCOMPAT��)����VWVAR �p��"�N���  �� d���Ң�_�DEFPROG �%�%MAN�UTENTI��INCEAUTO{�~��ISPLAY#���INST_M�SK  � ~кINUSER��ִLCK(��QU?ICKMENL�ִoSCREk��~*�tpscִ�(����Ɋ���_��S�T���RACE_�CFG ��jL�Ϡ	��
?��~��HNL 2�L��S� y�?�Q� c�u߇ߙ߽߫�����ITEM 2�+۟ �%$� � =<�B�T�\� G !b�j�v�&� ����4����j� ����i������� ��@�0�B�T�n�x��� ��Hn���� ,�P�"4�@ ���d��� L�p�K/�f/� �/�/ /�/$/v/�/Z/ ?~/*?P?b?�/n?�/ �/?�?2?�?OOz? :O�?�?�?FO^O�?�O �O.O�OROdO-_�OH_ �Ol_~_�O�___�_ <_�_`_o2o�_�_�_ �_�_�_joo�o�o�o \o�o�o�o�ot ���4FX� *��N�`��l��� Ï�ޏB���x�*� ���w�ҏ������ȟ ڟ>��b�t��� ��� V�|���򟲯�(�:� ��֯p�0�B���N�ʯ ܯ�� ���$����Z���~���Y���S���|��^��  ���^� ѵ���
 ��������d�R_�GRP 1���� 	 @�� L�^�H�~�lߢߐ����ޠ���������%�x�I�4�?�  d� v�`��������� �����8�&�\�J���`n���������	,���� )�SCB 2�z� O�L^ p������d��X_SCREEN� 1�7�
 �}�ipnl/g?en.htm�<�N`r�&�P�anel setup�}������/"/ ��Z/ l/~/�/�/�/+/�/O/ �/? ?2?D?V?�/�/ �?�?�?�?�?�?]?�? �?.O@OROdOvO�O�? �O#O�O�O�O__*_ �O�O`_r_�_�_�_�_ 1___U_oo&o8oJo \o�_�o�_�o�o�o�o��o�ouo�UALR�M_MSG ?7���� _zQ c������� ��6�)�Z�M�~�2u�SEV  @}i��0rEt��z������A��   B������7��%� 7�I�[�m���������ǟ՗��1��Ƌ �?�4����A��*SYSTEM*&��V8.1079 �G�1/30/2013 A 7���5�"�UI_ME�NHIS_T �  8 $q�T__HEAD��}�ENTRY ���$DUMMY2�  ��3�� � j�OUSEt����$ACTIO�N��$BUTT�ˤROW͢COL{UṂTIME���$RESERV�ED��j�PAN�EDATt� �� $PAGEU�RL }$F�RA�)$H�ELP�PA'�TER1+�<���H����H�4F�5F�6F�7�F�8+�INB�VAx ���	�STAT*�⥥1r����� �j�USRVIE�Wt� <Ġn�Uz!��NFIG���FOCUS��PR�IM!�m�����T�RIPL*�m�U�NDO_t�t� � $4�ENB~��$WARNJ��e���R_INF�Ot�y��_PR�OG %$T�ASK_I��t�O/SIDX��R��`�TOOLt�� 4 $X���$����Z��ߡ$eP��R�°�NU�$9`�U&�t���������E��`�OFF���u� D{���O?� 1��)�Q����GUN_WIDTH  ���K�_SUB��  
`�RT���t�	��$D�����ORN��RAUXz��T��ENAB-����VCCM���~ 
$VISʠ�_TYPɳC(�RA��PORTХ�A��C���N(�%$E�X��_��$��_(F�P��P� A��a��LU �$OUT�PUT_BM��ր��MR_���h ����+��DRIV����SE�T_VTC���B�UG_CODɴM�Y_UBYȴ6�	 ����ʠE��,���:��f�x�O�HANDE1Y��E�8pULX�P���AL_���GD_SPACIN���RGT�������0�����U�RE�����U��w�������o  ��RG��#PNT���R����� dġXr�FL�A���	T�AXSl���SW��_A���y���S��O�BA���zy�	$E��U�E���y�Ҁ��HK��� �
�MA�XvER��MEAN�	WOR��z���MRCV�� ���ORG9pT_C�&P )�
REF���-�i ��яN�b �b1��_RC ���� 8���M����M���� ��P�űG]����?$GROUP����<:&�� ��w2p CREǰ\w��$�Ab"vN!HK��SULT�{��COVE�����a NT6� �%���&���&ձ�#m L6��%F��%���'ձ����9�0� &z#PAu� �z#CACHO�LO V*4@1��E9����C_LIMIf3F�Rn8TDn8�$H�O��=�.0COM8������OBO�8(�� �!$IN_VPx�����2_SZ3�#2�56�#�512���8R��:TKQ�8o0�8�WA5MPBJFA�Io0G�?0AD<rIU�IMRE $�Bo_SIZ/$PM���ND� P�ASYN�BUFP�VRTD��E�D�A�3OLE_�2D_��EW�PMC��TUq�@0Q� ޴EECCU��VEM��)54Ro6 ��$���� CKLA�Sv�	�VLEX�E5G��� ��z!O�FLDd�DE�CFI�@�W� �W��<;�s� (��ߎ޵��QǠ�� ��_��L�#��8� hP �1��!���K�$��$=�E*�!}�C�U%$"eA7
�@PSKt4�M:&�e  ���TRbUt� $.p TIT-��A0�=�OPɤ�VS�HIF:�``��|!#����URO�d _R�@�+tH�C =u��L�^�p�o0���q�i �ҏsTI�!�tSCO'r�sC����S� ��SwS£vS°wS�x����Ꞣ��s�EqD���w�  �SM7�A���$gADJ�`K��UA�_{"u�A��g}�L�IN.����ZAB�C�����
~
��ZMPCF��G  C��J���LN�`�a��I��ԇ ���1� ��C�MCM��C�3CA�RT_6��Pa �$JT�N�D �1Z�k�d���p�����UXW����UXE�񞖙�_���u���`������ɖ��ZP5A��r�������Y���Dc� y�2v�/�IGH���h?(�p ���$  Ǡ �d7ۀ$Bm KK�]a_�b�#u��RVn0F��cOVC��O�D��$�`��Ǳǡ
�Iݣ�5D��TRACEW�V|a��SPHER�� ! ,p 1�G�vY��$�DEFx¿?%���c���^�(%� ހx���t�����ѿ�� �����*�O�:�sϰ^ϗϢ�T�IN�� K c��Ϧ�_T`�H��1 c���(�� ��(/SOFT͡�/GEN��K?c�urrent=m�enupage,153,1��T�fߜxߊ߀� �.�962A����������߿�36��Z�l�~� ������������ ���7�I�[�m����  ������������� 3EWi{��.�����'� �ѶSew�� �����//+/ �O/a/s/�/�/�/8/ J/�/�/??'?9?�/ ]?o?�?�?�?�?F?�? �?�?O#O5O�?�?kO }O�O�O�O�OTO�O�O __1_C_.@y_�_ �_�_�_�_�O�_	oo -o?oQo�_uo�o�o�o �o�o�opo); M_�o����� �l��%�7�I�[� m��������Ǐُ� z��!�3�E�W�i�T_ f_����ß՟����� �/�A�S�e�w���� ����ѯ������+� =�O�a�s�������� Ϳ߿�ϒ�'�9�K� ]�oρϓ�"Ϸ����� ����ߠ�5�G�Y�k� }ߏ�z����������� ��"�C�U�g�y�� ��,�>�������	�� -���Q�c�u������� :�������)�� ��_q����H ��%7�[�m��������$UI_PANE�DATA 1�����?  	�}�/` /2/D/V/h/ )j/ �/�$��/�/�/�/? ?z/7??[?m?T?�? x?�?�?�?�?�?O�?�3OEO,OiOvI� ���B�/�O�O�O�O �O _SO$_�/6_Z_l_ ~_�_�_�__�_�_�_ �_o2ooVo=ozo�o so�o�o�o�o�o
}L+v�H_M_q� ���o�>_��� %�7�I��m��f��� ��Ǐُ�����!�� E�W�>�{�b�����$ 6�����/�A��� e����������ѯ� ��\�� �=�$�a�s� Z���~���Ϳ���ؿ �'��KϾ�П�ϓ� �Ϸ�����.���߄� 5�G�Y�k�}ߏ��ϳ� �����������1�C� *�g�N������� ��X�j�(�-�?�Q�c� u������������� )��M_F� j������ %7[B�� �����/!/t E/��i/{/�/�/�/�/ �/</�/�/??A?S? :?w?^?�?�?�?�?�? �?O�?+O��aOsO �O�O�O�OO�O�Od/ _'_9_K_]_o_�O�_ z_�_�_�_�_�_o#o 
oGo.oko}odo�o�o�o8OJO}��o!3EWi)�o�U }������{ 8��\�C�U���y��� ��ڏ�ӏ���4�F��-�j�v�TCNK�$U�I_POSTYP�E  TE?� 	 v�͟���QUICKME/N  ����П���RESTORE� 1TE?  �]�G�A�S�w�mr������� ѯ㯆���+�=�O� �s���������f�ȿ ڿ�^�'�9�K�]�o� ϓϥϷ������ϐ� �#�5�G�Y��f�x� �������������� 1�C�U�g�y���� ������ߚ����� :�c�u�������N��� ������;M_ q�.����&� %7�[m ���X���/�!/ۗSCRE�?��u1s]c<�u2\$3\$U4\$5\$6\$7\$y8\!��USER> dC/U"T= ^#ksf#��$4�$5�$6�$7��$8�!��NDO_?CFG ���`��a��PDATE ��)�No�neޒ� _INF�O 1�&Q0��0%'/l?x8Z?�?~?�? �?�?�?O�?+OOOO aODO�O�OzO�OԜ>1�OFFSET ��OS5��_ _0_B_o_f_x_�_�_ �_�O�_�_�_o5o,o >okoboto�o�[ ��m�
�o�o�HUFRA_ME  �d6�;1RTOL_AB�RT932rENB�;,xGRP 1	�0���Cz  A��s�q�a�������v��*z�U�[x1J{MSK  �^uQ3LyNq%�I:%�o��ݒVCC�M_PAp 
�<%~VS?CAM1 *ߏ�V�����5�����MRwr2��Ҁ�$?��	с��	ֆ�Z��1B��5�A@��pp�pȣ� �o����������<������uA����T�Z� B���o�Z�s��� ��۟����ܯǯ �� $��!�Z���;���{����ƿy������ISIONTMOU:p�^�˅���"�f`��f`��@�q FR:�\�\0A\� �� MCT��LOGa�   7UD1T�EX�ϰ��' B@ �������ϙ������ �  �=	 1- �n6  -�� �t�����,x ֌�_�=���h�����z�TRACIN��$�4��� (��h��ݧ��� �������"�4�j�X�n�|�����﯆L�EXE<��11�-80��MPHASOE  &53k�޲�R 2�
 ��]�o������p�a������ ����� $6*1l������?������� s����������G	no�pqrs�tuvw  Z�~���� ���./f</n `/r/��/�/�/�/�//h$/?H/&?L? ~/p?�?�?�?�?�?/ ? O2?$O6Oh?ZOlO�~O�O�OD�u=�3��?�O O__LO>_P_b_t_�_D��D	��BH
�O�_�O�_o 4_&o8oJo\onoH�@�~		�3�
�
��Æ�o�_�o �oo&8J|o��3�
�
gh?ijk�@\ ��o��o�o����&�8�ƃ��SHIFTMENU 1>�c�<��%�ϖ�&���t���ӏ����	� ���?��(�N���^� p��������ʟܟ� ;��$�q�H�Z���~��T��[�K��	�VSFT1���~VSCAM�5ذ?��!�@`��^G�  A�ٰ8ٰٰ��p*�$���"�!�����L�̦MEP �a�/�[ T�MO����zR�WAITDINEND � �w�>��OK  Oյ���ԿS迻�TIM.����G��5� ǿX��8��8�%Ϲ�RELE9�h�s����TM��s����_ACTIV��1ѹ��_DATA �[�2�%��h�,��R�DISg����$�ZABC_GRPW 1۩I�,�q�p�2p�t�ZMPCF_G 1�v�I�a0�������MP��a۩/��'����'�s�8�����_����?������� ��/����V�������`�[�������� �����Ѕ������P_CYLIND�ER 2�� �Н� ,(  *m~��j���� ��%g H�lSe��� ��-/��D/+/�h/O/��/�/��=�29 ۧ4� ���/ <�~�3??W?e:�/��?�7��1A�;S�PHERE 2!M�/�?R/�?O�? 8O�/�?nO�O��OCO )O�O�O�O�OWO4_F_ �O�O|_�O�_�_�_�_`_�_oo��ZZ�� ���