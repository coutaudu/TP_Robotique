��   ��A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ��	��BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DNSS* 8� 7 ABLED�? $IFACE�_NUM? $D�BG_LEVEL��OM_NAME� !� FTP�_CTRL. =@� LOG_8	��CMO>$DN�LD_FILTE�R�SUBDIR�CAP���HOv��NT. 4� �H�9ADDRT�YP� A H� NGcTHOG�m�z �+LS/ D �$ROBOTI<G BPEER�� �MASK@MRUv~OMGDEVK�%RCM+ � $�� ���QSIZNTIM�$STATU�S_�?MAIL�SERV�LAN}T� =$LIN��=$CLU��f=�$TOcQ$CC�5&FR5&ALAR��B�TP�\#V{ARd(�RDM*}� $DIS�=� TCPIo/ }3 $ARP��)_IPFOW_x��F_IN{FA~LASS��HO_� INF�Oz"TELs �P~���� W�ORD  $oACCE� LV���OU wORT� �ICEUS� 0   �$��#  ����r1��
��
g0VIRTUALo?�1'|0 �5
���F�����4�5A��� �=��!y1�O���$ETH_?FLTR  �6�3W �������!�K�� �=2K�"oSHAR� 1�9  P O�O�4�O�O�O_�O*_�O N__Z_5_�_�_k_�_ �_�_�_o�_8o�_o no1o�oUo�oyo�o�o �o�o4�oX| ?u������ ��*��S�x�;��� _�����䏧��ˏݏ >��b�%���I���m� ������ǟ(��L� �E���q���i�ʯG�z _LIST 1}1Mx!1.��0ӯ���1����255.M����	��5�2
����0�B�T�f�x�3����� ����̿޿x�4���@q� �2�D�V�x�5rπ����Ϫϼ���x�6 ���a��"�4�F� ���1�K��}0?� Q����=��1�C��g�y��^������Q����� ���9�K�]�o�.����������J$� �>�$�%� �=��5�5�	1��9�@@H!�� X��rj�3_tpd���1 |�0y1!KC�0�m	���6�!�CP0����!�CONn03n�zsmon�