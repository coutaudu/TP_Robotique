��   ?3�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����MN_MCR_�TABLE  � � $MAC�RO_NAME �%$PROG�@EPT_IND�EX  $O�PEN_IDaA�SSIGN_TY�PD  qk$�MON_NO}PREV_SUBy �a $USER_�WORK���_L�� MS�DUMM�Y10   �&SOP_T � � $�E�MGO��REwSET�MOT|��HOLl��1z2�STAR �PDI8G9GA�GBGC�TPD�S�REL�&U�� �� �ES�T���SFSP�C���C�LC�NB��S)�*$8*$3%)4%)5�%)6%)7%)S�PONSTRz�"D� � �$$CLr  ? ����!������ VIRT�UAL�/�!;LDUIMT  ��?����$?MAXDRI� ��e5
�$.1 �%� � �d%Open ?hand 1�����% a?�? �" � �!�# �%CloseQ?d?�?��?�9�7RelaAx�?�?)OOO�9�6L82QO2O�OVO�3 @�?�O�O
_�O�4O �O�Ol__�6�Fh_@�_d_�_�[�3���_ o�_:o�_�_poomo �oUogo�o�o �o�o 6H3l-�Q �u����2�� �h����;�M���ԏ ��������.�ݏR�d� �%���I���m���� ���*�ٟ�`���� 3�E���̯��𯟯�� &�կJ����E���A� ��e�w�쿛�Ͽ�ѿ �X��|�+�=ϲ�a� ���ϗϩ����B��� �x�'�u߮�]�o��� ������>�P�;�t� #�5��Y���}���� ���:�����p���� C�U������� ���� 6��Zl-�Q �u����2� �h�;M�� ����./�R// /M/�/I/�/m//�/ �/?�/�/?`??�? 3?E?�?i?�?�?�?�? &O�?JO�?O�O/O}O �OeOwO�O�O_�O�O F_X_C_|_+_=_�_a_ �_�_�_�_o�_Bo�_ oxo'o�oKo]o�o�o �o�o�o>�obt #5�Y�}�� ��:���p���� C�U�ʏ܏Ǐ ����� 6��Z�	��U���Q� Ɵu������� �ϟ� �h����;�M�¯q� �������.�ݯR�� ���7�����m���� ���ǿٿN�`�Kτ� 3�EϺ�i��ύϟ��� &���J���߀�/ߤ� S�eߟ��ߛ����� F���j�|�+�=��a� �������	�B��� �x�'���K�]����� ������>��b #]�Y�}� �(��#p� CU�y� /�� 6/�Z/	//�/?/�/ �/u/�/�/�/ ?�/�/ V?h?S?�?;?M?�?q? �?�?�?�?.O�?ROO O�O7O�O[OmO�O�O �O_�O�ON_�Or_�_ 3_E_�_i_�_�_�_o �_oJo�_o�o/o�o Soeo�o�o�o�o�o F�oj+e�a �����0��� +�x�'���K�]�ҏ�� �����ɏ>��b�� #���G���Ο}���� ��(�ן�^�p�[��� C�U�ʯy����� 6��Z�	����?��� c�u������� �Ͽ� V��zό�;�M���q� �ϕϧ�����R����
Send E�ventU�5�SENDEVNT��z3�i��%	}��Data�ߘ�DA�TA��3���%~}�SysVar�SYSVY�3�>1�%Get�߂�OGET�����%Reques?t Menu����REQMENU!�2���?߀�;ߤ�_� �����������F ��j+�O�� ���0��f xc�K]��� ���>/�b//#/ �/G/�/k/}/�/?�/ (?�/�/^??�?�?C? U?�?y?�?�?�?$O�? !OZO	OO�O?O�OcO uO�O�O�O _�O�OV_ _z_)_;_u_�_q_�_ �_�_o�_@o�_o;o �o7o�o[omo�o�o �o�oN�or!3 �W������ 8���n���k���S� e�ڏ����������F� ��j��+���O�ğs� �������0�ߟ�f� �����K�]�ү���� ����,�ۯ)�b��#� ��G���k�}���� (�׿�^�ς�1�C� }���y��ϝϯ�$��� H���	�Cߐ�?ߴ�c��u��$MACRO�_MAX:����_��Ж���SOPENBL ?���������r�r�A���PD�IMSK�����Y�SUc�u�TP�DSBEX  -�q�U����n� ���