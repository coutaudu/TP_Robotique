��   j�A��*SYST�EM*��V8.1�079 1/3�0/2013 �A   ����DRYRUN_�T   � �$'ENB  �$NUM_POkRTA ESU@�$STATE }P TCOL_���PMPMCmGR�P_MASKZE�� OTIONNLOG_INFON�iAVcFLTR�_EMPTYd ?$PROD__ L ��ESTOP_D�SBLAPOW_�RECOVAOP�R�SAW_� G� %$INI�T	 &J_ � 4 $TY�PENFST_IcDX�@_ICI�  �MIX_�BG-1
_NsAMc MODc�_USd�IFY�_TI� gM�KR-  �$LINc  = �_SIZ�g�� [. , $USE_FL�C ���i�SIAMA�Q�QB&'oSCAN�AXC+�INC*I��_COUNrRO��O!_TMR_VA�g�h>�i  �'` ��B��!n�+WAR�$miHp!k#N@CH���$$CLAS�S  ���� 1��5��50VIRTU� ?00'/ �>55���*����w8?0'1~5��%'1�?���?�?X��O5I1Z;� O'O9OKO]OoO�O�O �O�O�O�O�O�O_#_�5_�?+ W?>5=d1 ��t_��_�_  �1~0��_ k 1Z; #4%B_�_��{1�1 �_%ooIo[o:oo�o po�o�o�o�o�o�o!  W6�1�S��Z=�9~0�� �r~1�tX{1>1~0�>� ���*�<�N�`�r� ����������~6�1�q �1� ��$�6�H�Z� l�~�������Ɵ؟$4�v6�S�1Z9 �)�;�M�_� q���������˯ݯ� �Ό�4�F�X�j�|� ������Ŀֿ���� �0�B�T�f�xϊϜ� ������������%� >�P�b�t߆ߘߪ߼� ��������!�3�L� ^�p��������� �� ��$�/�H�Z�l� ~���������������  2=�Vhz� ������
 .9Kdv��� ����//*/</ �6